XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�K�i���{�o2M#�K�C}�ž�r/�B��t$�?8�S_ /�*�I��<�!�61ֱO��8H��g/#*㻹�n���}�Iؽ7ewx!���|A�uh��nl �U�Q~Ġ�>%R����i��5��)�z���E!/�/9��ք&{��? ����1��	�lb��%�g��~��ጆɪ�"$�@6������e���MM_V�@M��6X���Ӽ���0�4ԿR! ��}4�(�y�ģ*��C��*~@�݅R�0{�i}m�%��6s�-,v�C�X1��\�UӞ��%���;���C!v��*��O �^]���5�8O�^N���5p�UnW�MVJw�������ĩ3 _Cq��ژ�%�T���_n���X�}���A!g���Y�u>�R�W.��t�bXnJ�K*D�n��^����ǒX����x���+9��&9!l
�ˈ���Ψ�CI��N8�!�y��x�e%SC�(�O9*9�u:F./�AŴ��yϟ{1�Yu�����?ҿ�cn��[a=a>/��ӌ�yt!�&���׷����	5���rT�cf�}ｇ�_q���V���´��q�Ԫ7�aC%����]paEdVֵ�W��̄	��vA`��,FD ֌�2�n6�~[28�؊��:C��@Rx:@�Ҝ��ޏzxT�(�Z���&x?�s��z���Ṝ�Klez�	@�m-1A')D�9AǍ�����S�Kډ�끦�:%R��G�XlxVHYEB    9de1    1670gd�T�3���� ҴӮ՟�f/U�>_� >M��bz����i�{)6*�@}y��B�~jI�2��9ٟ���$��'�!Wj���Q���M5�<˪|L���<�=���r�&&=L�p�X"�N٪BYD�LQY�k�Y%Z��J]���)���F�:[�O%�GM'��)��O��$��}a��D��>�I�8Ȅ����qI�"��٢M��ܠ�"�7�׊��+ p�@��[�2��v-����l�SIP%�p��WB-�c��z#�Fǧ7�L'����u���#���!'�d�H8�*�v�����Tzg��ͽ87~��uM��/��o�0��)��^BrY�q���m�qlS|��}�t1�0�^u�)��
���UL�4g�̬��Թ�z�H&���*�q�0�~Aϙ�mA����?S.
a' \]�58J�)��iE��X�J%R�=Co���w~�ɴ$����<���j�ú`*}�/�ŗ�?�^`���L*���~0H��ŏ������|��7�*V����C�}ѷ{�����"��Ǒ>n\H`���}#��M&�e�?U�;	�CPDj���������}�ŵ��/8�8\{Ü�	-�{:(�m�Q����^�p�M�R��KH�
�gZk�N�w���0#1�a��LxR%c���\j��� ��ӗk���\D�K6r<�\\��
����	�� <zfJE0]�v�*�"s�j�66Ց�ު��WF���@#&�4���s~���s(��K�9�6�D^/��uh��*�
���+����SՓ}<��^|�*.���]�%���['!�7n"����!��L 6:�������W����h^J!���L<�|�Hv%�t�{r��\���\�Y��N_�K��[�#���K��NDn��?�*K��|�=�S���`36�=��A��h���R��.\���^� ��|�>����C˻k��qwR)ˊ�׬k�*����E�5�Dڄ��Z�~���1��9 ��{�6���Vl��������	ؘ�.�a��] �oRX�9�E#�.ܾ������������]�RfF������L�z���R�ҍ������n����u���^2S�E(��n��	�]�I�a&e�~�ָ�,[���igQ:v����"�Q����~�a��*/XG/2<�E%F[��ȟ_�Q���q.�ה�
eme�_� �_����4�kb��(1�otj��6E�����X /B~Θ���. �\q�T�4��Ltۆr�d�*1ڿ���r8�8%=faQr���y�C����/�����x�d��e�ރ��$��3m�+�	v�`"{ٱI�l���Rn�#%E���ր��s�mғ}$=�ˎj��=}1.z��~�L�ϊw��n��;Ŷ�:�=X6P�1�ς�ec��u]s&����R�;��6>څǴ&��m_��Jf��)m2<<�-����xp�G��NN�#'~c��9��܇���`h7@��ŭc~�h����/3Za���S<�_W�A�׵�.���sR�qhy�삐¡!)���$`x��&��߾f��\12��G��Y�1��~ِ����|���^��ɫ|.�Xv1��̜{6 $O��&�U�� bW3���*G�A��+���-�s�����#�.�*�|���+N�M�q��=�1 ����7�6;�zκ����8��A�M8�� �t�����,�ǫd�M�M��H����N;����̖`�1Ԡ(�ˎ<�^����d���5B�˶���Γr&'e S�+�!���ǴZ�Oq%�
B�#�`�Q���ט�e���f}BO��d�Z�2�+�^��s���`KS~u̷-,�#�^`�9k!�N���|PH��T��9��#���T�:�	�PN�^uO�4<	��M�0��*F,4���n���3�&Z��^�������&|}.��g��42z}���d_��։M���~����hSu6�e�b��i�����V�<�R8@�6��+js�;)�l̲���<lR]��6X�R7��_�dV�9Sdx�/(}(H����d�'�\?a�w��+ԺqW��H�a�`5]
�,<�����=dP����+}�+��@��ҏt�Nn���5��j�)���x:r�(�
�PDn�x<�G슢z`�/a�>8�U�(��pE�Ow�Y[05p4o���k�T�WF�nc��(�MWDa�1�$V^�p�g�� x�	vL��B}>&��9~�q��s���=��}�~��}��Kx��;�ä^s��k�q���Z�����������q
��u�Ҁw��A<LrHjZ�F9�g����VN=bŤ=�ʄ����ѢϾ��J_���<�`l����벟gJQ���V� �k���g�Z�C�Ls������C{9	bcW�פ�7ý�mJ����^�Uy����e�0c�,��yP�-rz�����_�ea��$�J �h�ߧ�����Õ�34�:��w|d����L���\����c���1����L������ɲ%�4Y~�A�<f留�'���B�Ɇ�Ō~<E}��51���ш�]�*0��T'���w�3�����4 �ڃϱ����d����k��1�uš�<1#�$*ȅ�s�Q��O���3�]3t�I���9�;Ρ��C>k�9��\�7�m*�K�v8(܂�	l�fR��e� G�'1�cݽ�M(�a˂	q�7�{���K�p)����U�*�v �9$d���a�_O��lf�t�y����X����h~�fQKwfk�řŀ	+�'&UYC�X��h*���W��ƀ�#�ɐlo����[�H�]��YA�E��5���"�PǿWt�S��8��Gv�h�E�,����{O$�20P0_]n�\" �N@C�4�[��Ń����C���Df����Bt��Fɷ���9nJ�?����L�q�_��D�E{�`Ł%Ih1�{�C�J/%���<B�L�=�:8~ ��~����ڹ��vj�������u���Q�S׮X��U{"���ԍ�/g1��񎖓Y�>2��]:$�{-���q��pM�Z�';o��!u���lE]N��e�xI¼�[j.��5��V
��_�Wl�א�Q)X�R�(?̪OyAy�f�G:3IJ�'���c�9O�J��8�������9�,|l�+�}=��~��Z�f?�缙4��T����c��p��N�^ ��Ğ�<b��,1��qm�>k�l̊��w�X<����﷖��(n�6[�25��9�`d-ǘ5����6W�&~h<yC#(�g�^V�������R�)�-�0����{����`0{���U���j���������\Ӝ��7��~���!����TZ�>�8�5���<��qע�7b�%�H=�{l�{"��:s��k j��翩���X0��-A�y~�;�bv�Pa����u�q�� ��BYg���*cFp�E=�<m��j�F��݋No��*Ž��S�}��/Z������̘��� ��g��ݸ_.��XC�%�H{3�&Ҝ2�=��F��^�Z�#H�̱��zE�fFÇ���Q����LT�_�#��E
�����|0��'q��������0QD#�B��%MF�#�`q�f�����7v%}A~��p��g�cW�D Rz���7�HlD���έ�F���R�ׁ�[�຾~����GU\�ǌ`Ojv׬�����/g*���eF���z��뜡��en�l�N�*ݎ(�����r[5h�ԙ�yZ�`�jB|�^i
:J_�!E-�z��dt�gd?<�~a1<�|�:�b�7E3���o��S��s�/w}XÑ%�xZ����w��Yp���)��\���頋޴$�c�1Ѝ<d���.b�X�W0,7�i3�eRIӫ�j��&��K�V����y��Y���^vkw��q+ސm�.�j��9C�)��$YGI�J���Ӽ3�_��ԟ?������xk����
�j΢�<�y8�|������:���l����
$T���dn$�΄��;�e�#X���Ԓ>Ѫ�����;�ŀ�%{^UB����m(VA�U>�������k�m���3�{�����ha��S(�#K9qۮݝc��i�O>�����.E�a��@�����h�SK*��eS�ڐr�
rs�t\Euw�~�ޘ��Ob�~���fBƇI��E-�/��.����P��,H�ϊ��5B˳,*�u����Iz��#�o�Oc56��+�&E(��c��,.�n���e��BzC4s^���iѓ��d���Sy�S�!W	�Kp��׿� �E�����{�SL��z��.
w�2�+<�k�w~�;p�� �L�d������E1�6�88��1�ȃ�$�)W�N����#�q}���DQ�}�h/���(����o��@��'��>��i9���s�Y�(�K�grox����E$�U"Inث�x;��Dr]��ﯛ�TÌ�P�ڃ�=���e�X�r����
����T����}0�W���)K�C��M9�{�¼ؽ�J �0,���W�i'Î�m��hq��yM�ʲ
�_�]u�7��dii]+9mTB�~mЋ�H�&�?�����\��<�ζ����؎�ͬmEr��JKpxs3�Gў/� �ȇb�~�B �\�`���X!�o�GP\e������8$�Ģ��r,��B�j5�;�;k�F�rߧx;:A
7wz�2f�m �o;����U�HJ�pH>�
����,� ���F?�Б�j��TA)Q��+7�U'���_6��ek�8~sl�'e�&�oQ0f��V�(��nyģ����Du�B[t�K
� �
<(�m�VS��9ы%�_���t
���R@N��-(���_r n%;�A�����o���EΖ��S�I/O�^K�ҿ�	�z������r(��g����V^�z/m��^�כ�.[��ڿ�I�_JE��L��t�>BQ��?��M�dB
;�Z��@Ju��~�ر�={x�����
�O>p2$�������H��>��U�зW͇]������3ƨ*�fC�4�I	I� �Q	��z�ߏ���	�,�_�+c�
��:��a�9�3ς��W5Ʒ�^�Z�R��U����������jY� ��"�ت��@�+ë��>.B\w��iQ'��$�RJ�]ܙ~�M>���ad
���s�^�jM�nŞ���[qGc-YҷA�XZS����Р���O]\]$f)n5UmנJi4,��caæ|�V�l����	.�;��,����p�5y޵�tT0���v�U�I1��h.MȠ���U��)�y>%E틵��9�?��IXZ���ɗ3fӴ4>�O9�#���G:�<�<<��[�p�=ɹ���eA�橈�ej�<C�t�����I߲�c�W�V����M/�p�SC�dk�ĉ�~=� P��8gV!X�M�A8q�pD3-��ڬ`�v�Q7�"ѩD�hp0|��Q���*�;H���sľ��s��y���A����Cd'i�x49>�,?���<y�v��T�8� �E����wٍ�Ӻ\L#y���B;�,H;��ת���i��];�9��゛�)��~�N#1�7�� ��:#�R���>~d