XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������n���˦ �W��R]
ㄒ���V�ee��L���iZo���.�0�0y��{���|��8
t�kΜ�."z�a�+cj�Ԍ{�/�t��T��T �k��Q�[`k���#gpQ:o��l��*����{�PZa���|'�w U������r���1��@'�'�=�Hm�{�t��n�p�/	�������5�<I���RpUsB����h�s�3bP��@#��_W���]�is���\��n��N���#���Ru��枦V�'s�Jw-/��d���T��7�r�6�l{�T���R�A
�c���~~�c!2�v�mU�h���+�2Hˀ"� ��y�.��E�G�d�� �t؍{G+�$e׮�#�ر�I�R�O��Ӏ�Y�=KǒK��X&�����d ��Hs�\ǫ;�t��\�CGK���rx������rƤ�8�Ɗ�:�Yy�zO�;�9|;�N$a��32�Y�Z�7bb!	۷��/a�4��s�}��~��ຳ[�8�5����c�V(<��!? �W>���\~+��9[4��~���A@Ғ�*p�L�S��٠�я��a��Pz���͏�i����@�	*xQ��?M�d��ӹ��|L�[�����+� ���R�hZX�ܴ��p�?�!$.�]���Æ���Jlyi�FYQ���uûﲔ殍�)�1���҇�KX�N|���3�5��܆V�.������|xV{�~��F�wZ|�X������3XlxVHYEB    fa00    22600|Ϟ�5Aᕇ��]{�(�;���=��v�	�輄}\F���H��cL�*^��
f���<��l��*V�Flgxg(s���d8�K��)\OJA�<'+L�e��.P�7�ͽ�_t�>�ȗh�D*�OPWTYXo"��.w�0�f���W�����p��j*�a�����"�p���aD��a��1)�Y����� }G�7`�S�^��_��H��:t���<i�� ǧ&����:���S���K�V����UY2��^T�4 �&%�����࠲p���̺�۰�n��Z��{w����V��9
ԍ�-(k�{�rH�S¯�Y�a7_ф9��%�0�T<�g�i��]������"�J:�k�s�x�2�V!��m������A#�_:Iٰ9&�;@X���3�bB�H�8�Dk�߃sh٣w��ƺ2rB^� ���u��V�?*�G(&<St*��*Q �J@�v2�!m7�024�U�W-K���Q~�?=x�;�B�r3����]���?8�--�1#���H�5=��(
_�A@�.;udӵg�/���([��+����:��¤G��tR[�~�3��м*����*��G2QH�Sa�g��JrA=��zk�_\Af�Av� �P�����̫Z�Ŏ�t��_~e��f��&9Q���u ("�Q��8"����s�O���9fX���H\ W�G�{K��;S�
9�_u�E5�r::h\⚹�Lk���%#Hz���J�}�P}�C)g�������[}[ܽq,9��>4w$dn�>�R8�"�B�KB��IN�=[pw�MЂ���wb��^q��AM��#~��7��VɈ:�k�ED@R�i VS�e�`�Y�$�A�R*���&�zΰ��A�! U��zP."�b�2��vNY��ڍ����U�C��������,�w�[� ��$��x*}��+�a�!�|�+�n��	dӤ'Z��S��Jhj�tA��F�J(Tq��tJ��EQ�91��G�����-!�Q�ǜ�۔4|�p��XK���aK�8v�ϧ��m�DJ�L��]�Ќ;/r�>����W���0ĥKӒ�cU��Ůݬk�W�NM���o�4�'�>�Z5,t��-\�YZ����v��`|�?\g�PslA�K��l��p�I7��}�,%�0�����g�)_^*�m�%lIC�����Hf�7�x��O�s%w�����.���S��n�� �����c�%��4�2�S�6�ږ����@�0�IR8 �:Wq�.�De��"}-Ģ5ҁ�q�8�XS��,�����ـc���<��T}��-~�kX��g�>��
! ��GȊ"6��K�'TDca/+���P��9r��XI0Iݚ�%R�3���u���/<�"�OU�Yrty�i#��� @�o5nq���v:׫�59�~���x��ތ�\z؉uc*I�Z!�gF�z��A���d0�<���`�@�v1w�xjp��؝���o� �$�C+,Ru�#7��)����g	� ���v�8$�;��� |$'@k��x�uΉ^�5n�Aϰ�G���QlJ����8�AO��fNC�)�^2
�a�T�|���WfLq5�S&N��p��E@eɶE8E�;������SK�~�ϟ�+��~�D�S��[.gH(�RY'~�I�%!�jʉM�v�jb�nrB��Ε��ʶ����W]]7G����W�ZCl��ƫ��!!x�t�ZMOa��2~bG���6@}V�����B6d��YE^�P�7�\YkN� Q!���V"�C"��0)�%�ݜ���QK'�OM���s���nU~!j�f�����z-K����w/�P�¡1�&����h;5?%Q��_H9�=P)ʀ翃S$�m>>3��x�8ܯ@���4�`⫩q���@���m���o�O����?!*�+L��S�_,V�r��=|���tݦa�ŋE3݇z�C�4���P1N+�ۜVƧ �1��^��r4�������c��n���[��G˚��~�?d�^�T��S>@nȎk�[�S��+�د�B,�xI����6�YU[����'�c ��()��������X\x�:���_f��[ք�b��&�a~�
U��
�e��Y�ox�`#i�i��gI��������Lƭ�l�g�~�xa�N"�_٦x��o���0o�`�/�9`�2)L4�Sܢf���h-�n��0(�SPB���l�n��΂ע�^@����1-S�����}��yR�/�NOb��QqĪ��.4����DU���5�1BU��c�ƥÀ�Ud�f��� ����a���M��`r]&/�.�\,���q�^
y(O�՜ 繳�a�>�(U��$�(�'<�,SD��h��Q%��Aǡz�̗��'�?1��&�d_>��G���l������EZlp�(�������
"!�ٔT*�C\I���v#�17�>Ǎ&XB%c�q�iP�{C[�z�_޹�$�Ȕ-�X75u��OqR��6�H���J�t�@�(]���c���;����$��4�_k���������d�("��/tY�*{mqn �(�j��PO�s�����[\l˽1��yM�ۍC�U�,�G)+%N "�}�ڎ����F�⮌c�@ �t�5�����U�
� �-���)ɤ�@v��[yi��yG#��+^����?B���c�Ѯ��0~[�>��rbdJ!�K���E͡��� ��Pe�p�;��������a<V�{�����5�#��,���p��Gj�e��C���T��?#��kI�i��E��8Gq��'���|�����`yܞ�᰽�c�j,_��6k��GQh{�d�D���v�D����<�hH��H���� S�y����Gڦި����r�uh��ipl�F�S��l�&=���.U�����Ɋ
h�Ì�Q�ɢb��1�!�����jS�j]~�dl����{�s��x)~x��]� `s1Z���5Tڟ�E��Ac;���_�G�Ea�.�y�uH��>�~�cw�5�!e�bbC�n3A.M͵#�e�Mf��Ͼ���'�׻�0��ՓW�M���C(�/y�P J���aSZ�V�5�\�o��S��_��*pN;n�ݏ�m+G���RT�W��4�?R��(u�o�r���
� ���T��������YXDG.�Dm6|L�y�1>3�d��J���Z�>g��%�����*EC�4}��	'�#b��FA�V�M��}\!	��P�*�4�z�I��X�0�����;`��R�E�#Y�8[�#�j��`
�>����L�� �Fogp�0�Ȏ|�mϗEx��ҡ�c*���1��6�fH�%K����������d����l��٫}	9�4nf)B��֒���� ��qi$�����C�T��#V��f*5�P^"G��(�T�v7I������AZ�cO#Xs���w���^�b ��#���R�K�X�UYvI�����;�4�jD�C�,)6��3}1�D�T����ʤT����,���\��Y�|'�!	ÛoT-�&,�D���
�غL�6��Rx{�Ql��p�C�+ �̜e\1����Oq�g;�f\�{�6P���4�?�)5��f���_��eޤ�A/8��fж�y6j�g@�l`^�'
W�}x5���y�Rޢ�l�ՕQ{y�b��փ��Sd������{E���~�L�������t��l���\�fZt�L�U�z�W�F:�bUM�18d�[��}�����:�Wp�j�un�����kΣ)��>qX;�6�7�F�;(�t�t�X���B%��g�N���S�+#[)����I���M҈vy戵H�<�����P.;�p晗��E�B��|�N�����`3��A�U�k�y�<�.���X�]2�鯧���:�"��d�F�Ɏ�/r@G��i��e5��ҹK��/(?���؞8��=�S=C=���DC��]��˪Õ|�C}J&
�/�:n6� |Q�;|0����DjT�~�'����A�?���^m�5�SP����J_ ���_�E����4&W�F�������\�\.�E�ӳ�7-�~�q�����=/7��>���L����y�Sv��=�g,n�s�0�y�$��J���_^Ԫkvi���'tv�R㛓Au'n��u�ǉ`�^`B`pZay�g�d�Ƈ��U�<O�\���#��p��0}��51�v<�B)��H�B�����Y��h�>$��%�R��T�&q4�a��mT���a��`�McT��5���q�P[��>E��H��4���C�+<��p"��L2��@�S���_e@�"���-v�N�Ü')9Ꙗ'ȗ���,B m�{xtF�鰎7�+N ��5��h{��h���dL�}��"�����5�j)A���%RR���WyU��aɂQ��;R�)Ț#�H���P(�%�e	�(\-�Ӆ��+y!��� d ��M��Ճu-��Î����'�L��ΞM6�-����S�������G�����Q�w{c����@��n���)ߚ��y���R�|ېԷ�\b�Y�ז����Г�� ���,�q�E\��{X���������M�Q��$�U�EbZ藾E��~$h��v����o`F��鏉n?x�F"��(�֠������v�[e;��mA)^��u�Y�fv��4�q|�_ֺ��ґ2+�W�8g�9�Ͷ.�MDI*�:�i���Z&��+Ӫu�(n�a5��!8��Gݡ���(�H�ô/�	[��
n�M�����K���*թ�.>`�tg��VR������*��$e���^������ܒ����%f�϶���ץ����o,H�\��1�;����0*��+�I4N���w'�4WػG1u��?�^:���iF=J.ӽ���vjQ]�� ����A�M'���ar(_���hS��R��S4�Xt�湐�	`4�t-?a�cE�+!Q-�r���o�:�V.n�ȯS���|�!���W���P���U2�y������QS)]�e�e�ҕ�Nx�L�~�d䚅z� ��2ӟ�;��G��qB�[tpXI����?�~oɍvZ�0�w
c�y�XΧidk6���Yy�W�S�P��zVW���JUc���f��?e����w�����Ĳ��Q�i��,�$ǳIgU��1�����k䦱@�X��0K$$8Ob�e+='娑�KS^f[�!�J2'BM�Ƥu��MV;wK">1�c����8[iÃ��Z������ҙ��E�C��kɿAi}%���w�:�ȣKB�~-޳O�Z��FI���;�����8*Il߰���6��˭��R��u6a�X���w7%/�Ϲm����J#���"_B��De-��]�w��L��:Ņ{z h��ԖDHq/n���O��a�������YB3�џr����3,u:|ZG왗z9��,�Yk��{s�%����a�J�MxAf�`}��8(����
\F�S%�s䞨3��(֬� ��>����>tz�3�#&���330!��.~�]��I�`�D���1��Ah�k�f�q�)��Z�9�)e� �n �!�s��$���Q�l81�n�������RC���'%���ٺ3f�#��_�i��
�Ԝ:����k?\f�lf�J׆�P�L�2�����Pl��c*Qgc���iI�ݫSP�X
�� �L���6tCEs�!R�E�>H	"z욵�X��L"��ǟI_�Y/��ȧR��G�X��V�c�>�c��CI��&뀣}@�,�C�ʧ[��7L��6�m���D�&��+�\�.Z�S���9@0��A��&n�7��v���|2����z̇���ٛʡ�>����If� L��Dr���AL=.*@u���[���Q],n�i@#�2�{!��Dt10���I��)�0 �t��5����3]N�0b޽�`�{�,Z  �1��a[����j�0y@g}r�<��JmyG�E8c#ۑ e��}�ַ�qx�mez�M��w,J`�8��l�9���3��R���4�4�(,0�Iי�^��)���Zz7��M,ɐ[�	yo :++x}���3*���Чp����R�����\�Pw� j� #0@T@�D�7�S�N��?������Ab"��h5���?��n%��}W�
c������V�V��'�M�]�2����k��!*~���}���W�v F��_'��G��+n��US��-�n~��ͥ� �Lo��Mn�zp{�^V��x��uߙY�Ԍ�/(Iyc�އ+ J%^��M�q���m�ƈQX�&l,t
��C�c��_��]`zh�8�����i��	�Z�L2ț�caV����ūa!%4�Ǎ�]22//�=j���{��?��K_\��h���ﺰŅ$�>�WT��aU���>s��&�fh�Ng��?۔��.��s���CydGGx�V@���Z[DFZo<�l�c���0C�ni�ʒ�����	��F�b�mމ��!�V�I�;!�"9j�d�-+m�飬X�=�$���_[�n:�����h�$KNS����u��k�������z7�8��wwڃ;;hP�(0oNhM�>��[IX@�}�`(cm��,��#�t�1@PuK�N���\���B�
��d��MĻ��Wf�U���o�����%;�A���g~9A���J���^�ȪP����h�Eb�N�ph�SI�0؆7�5Ӊ� �} Ϩ YBv�`��*��1)Ȼ���+��9_S�_�v\�X}G�0�)�}p�?��j��j��×/h�����1�U�*1���C>�l��ඏ{�؂�D��#}�˕�n�oܨj\i(����n��2��<��ÞmhXP[�R�abS��)SQ(~x��Q�!p�*�!j�#8�t�.�W1�o����}���'m02K����l��@{s�9��M,5����K�f�}�=s��Y#��,�!�Q,�f�\��B�o�|l\�T��^$�q�4"�K�S���S�m�s���%Ӗd�B	���r�;�Q�-Sx9�*K�9��bkp]2��Q��!{1�������.rS@��Fz���[���t�����W�~(�a�䏖��NItR���X��O� {4��7�+&���P����>,�3'�`0��|�-����P���ୖ��#%��ހ���Q�*����R.Lz����>��_}�� ���k~c��s�IT3�ɳ#.͝��o��E��L~�m�{;��i��sa|7��prea%NO[���:E�O%]��iL�C������Q��d��GXb/N�����yǏ_0\Z)	�_�����Q
�7��m�n�f�xت� &f�d�e}l��P>u&�G�*O���&��a�Jw�E���D�MIg.�_zq$�q�T* #�"{}�=|��(s�m["UE�)�gr���k�
�	���lg����mS���&�A-K/m��~Z�a�)~�:q��,P���$8&����~�D..���Ǣr.W8�Ϥ��5mf����������3���3ʮӅW���ɨ(��d_S_R7�3�DL4ܕ++��V�"J��q�蘔��	�.�����nr���
���L�e>�V~�e(#ch���d|�׷��T�A BQ0��_�}-���O��9������N0��b3�p`�ż�e,x��#�4{����JHiH��$�Y��ί�5g��S�e.9Z)��: 2o^V2 C���JKT0/i�_]�Ϩ�Nԭ��h�����k��u#9�!�Y���\�Ri�������Ǥ4��U^Ӫ��A	��-|N��Gb�4����s�l���]�^s��cX�(�H	T6�	��j�'6����W��� �o8a�f�g</���E�فR*z|��L�J�/l�i����>5�t��4�0��|ʷ��4��h��^���g��ʇOw�����PϵKpV¡�UdK�V#o����cq�.���ց���U�C���J�Qf7�?�y0��k�?��V�]Q�>m�(F�3.�K����d@2>�M�6�<��e=��>S�>�G�GʛU7~�S�:J:鴲�y�ʻI rTXo��F=e
Yi���˭�c/5�}�<�#~w0
L�����Rsh���Џ'��Ap.����W�� ��o������ܦ!���gK�V��K��7��x��0��,��ih&�2@!x~���)W*mbR��a���My^��춇����i�����wTVu3?��/_0D�
S@e�8@O��)��O�?{����ܓ����x��#�
$br��x�ua�\��]!�(�V'�LW�'\eb���g�b������9g#�#=�$[5.��%�JR}�j�D� &���m�n�9�r�,1��(�m�PQW��Q�'w�d�A�asw,q�d��i�d<^�Ybh_8�2U� �J7qR�Qq�q�y����&��f�ތ��-��JM�AG5��M�&���A;Y�n}B(�
���@~7#���9梪;"t��B�S+�:�Fm���|�I_�U����^3�hU�`�����O���P��-�q(���#�([.�8���1���ܢ��֑u��!��Q=P�6$�%��W���0��9�U�ԼU~`VG�,r2R��XlxVHYEB    674c     5c0�����#��B3���R�%�A���L��"���k�և0 /%47�Y�A9�8��^,EOe�w�m��5a&8�Z�{���u��"B&� 3����Ѻ����E�Eg=`�6���Z�E�Z�G�	�����#D����>��׆��-VeI^�{Ɂ�3B]�
!��(�J����+�y�%��L�Tw_�����>l����7i��
�c��u!�wbP�lE���xiϖ��K2[�EA ����x@�������,p�q�.�v��W��{QU�I杀�3K ̓�G��tY�^��&�5X}0�*fo�-��K�5���:l!���v�e+�D�����Y |�蠽�˕+���yCH�ԥ%�/��e�`!�P41��X������H��ID�	l���ºAG��x)��ؑ'.��kvJ�e.xkɒG�gm��U\���W��@׿Ɠ:�%e�_�_]��le��DG�j�x�ue���Xݕ5��&0/͚�,"��B-#����y�;'D�9��Ѕw�EG5-���F�D{�}�VLs�3�~�'�cGrRͧ��X����b�S[.7�`��V��U<�\囟n9��h���U�ځ�ޗ2N+����=�xf+�[ʺ����L�� �[_6T�t�먷r=Ϡ�-�7�zJ���̨޶���*+8*���];��#r� ��y�f�z�z	}j�s4��P'W���������d���p]����ѕ࿵���<������:���(d�*����6��CK�"(+0���R��#�z������b�	PQ��]ΤG��=����u��I��!\���];n�Hn~'��vlL���Kj?�oI��^¦��d��
G����X����J�pNY��B�~��dyvb��u�&n��{Xs��w��vsq�5ѿ_�=���_��u臹$���+v�ym��΀b�9�@����4�*��0oY�_@��Y�bHn����F)������n�U	�7�Z����#4�W� $�
��Ⲣ$���MC3�tF������ᯔ�P�u��x��Ӿ�^
31��v�����G�K舒ǡ[g��?N�b�� �F��/�?�ǹ����ب��	=��W�w���/��?P����@�_�B�9#PG&�V�H�l'�x�@�M�T��ghBz	9�$V�>��#�HEe�-�cJ��rD�"�&�x5������s��x�ad%_�5o��.��H�r	�wVq��R�*�[yP��V̭!S2������*��s���7�Q�'Iw?d�f��m+R����l9J�&���.��E��^@�"��o�!VܣBt��������!_o? ?���:Z� r���5���p��]�җuO��4���<Y��~#$.�fv�МJ�nI�6���������F��C(G7��R�4�g��6�;��%\�)pc�ň��q�>�xm�*jS�O�;�