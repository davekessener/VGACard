XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��#'��HI����>d8��.�Lʹ�X�S��������h�r  �1�ur��$���j�V:�!|�-��c9,g�.!E�9���o��'���Z(^CBS[IS*��ooE��=�������)�5���0���8v~ϷaBb@�ʸϒPO�<�	E�;�s�Ŋ̱���X�(S��v�!9h�s�?Qt�7c`�sAI�����9���e(A�(�=E'ݢ���C�WQ�$����Q�E�@0G8[��꾞�!��~�`O5q�M{�5FŚ�)���P^C�A{߁����%�D�wF�z�Gl�~�V�q�(:'��d���4,�b� |P�}�4���.ؖ���y�WZ�=�@W�G1uѳ�U��| l7	Ɔ`�[��d0l,e�xm�3���ڶ�p2c�7HZ�;�*��%�i���(j��6�����_3��O����ݾ�Zl�ʍVHP�3Y|1��v�%�_�iO����!��ukg�/z��P��~>�!z�*�/�p�����ju�Il����>X���p"�b2~�Δ�]JA0��S1QF#��O	G�Y���)+m��'�c����ޝ+�`j��Pr Y5�[�F�V��[mV"�uAiѭ}v~��۷�mB�djll��?6��#��9Y��g!��E��2������mg�9����.	CzB3���ȁS���gD�08�P�?�!��ŕ
c�|���c�(-��m�=W�H$c���$�?((�v�a�H�n��Ӄ�!`�4XlxVHYEB    2e55     b00:�ϋ��_�mvè���������h�2�lvv/�J(���b���ظ�>Գ+�x8T���<��̹5�x�`i|��AK>bxCM�|�c+��Q��r�>���G��j����#�+�ۢ��������:Aj��+�6|ŉ�ǭ��jkpYv ;��.�ne�l�D33�-�zũ~���C��f$� �F�<�ں��܆��j��{t^����"����tT��n���6����\|i`�~<j�Q䖴�zc�(�潃L��B���X	��Gh�W\>� ɲ.�D��󹴐�A�:�d��������~1��J�o�2e
(���mZyn�|�<�~�˫��е]��c�G��%��L�5��-M?<���n���gԌ�Agf:����k��w�ݞ
�X]8غ��H%��{h���y�h�Ov���`tv�+?�$K�P#ͅ\o�$�?��&��s�SIJ%R ���w��帋������$ׂ�l�����0��g	��,{����k@�Ƌݟ���≍��e�E���Bz�K�c�*������S�"B�����Z���T���%����]��U���۬�.h�~_)�1Ȳ�^�փv0��=�B ���,)ጱ�����=%�$Ŏ@zj#�v�
�9gXH�Pn���q����m�4��\�(����z4SX�ii�|5����Q�=�����������V��-���%Х��Ū{�K
K.*�TC��L/��b7a[�kx�B+�K�|� [��N��72�|ՙ�̯��������zF�n�Uv=6�Fn�4���e�|�_�	�G��r�VI�(}�e*�&Q}�P܅�E�"�̈����u����C<��~i0���b壆"ߚ��EQ&Ȫ!޾�%E���,�!}�~�u���L&���o/�c�  ��Y�y ���?U*��(���t�D>�sM�
qlϭE�Fy�E��`К]�R��sMq]�	&I7<|�H��M��w#;�$DVG�5c���I��]o��*�̴�a�\�(��jr�2�|[��P�g�����B����a̙�m!e���9�X�nǺhm�Y*m�ox���v4�����e�P,�r��?��ZdG���s[Xn+?�@I&UC\���l��/�?�ɋ�wl�	qZ�{�G�OO�6�n�q����_���	}�i%N�!��0���/�dd��(f\����ן�V��o��陫���Q���S���-b�C�'��`LyW8ϛ K���$��hzA�ύK`B�Nq���T�ǻ[ҁ}c~���씪�{��.I�β���Y�L{_	
�N��^)u+���D�����R~P���v���v��/uߍ4!U�	�ĸ��epRoR�ui�$��Mp�-ԙ����	�Vu�^��_�u3��A�6��=Nb���F~9z&�!n`;C�$Xe\ϓ�/Q0�5��ޗVZ�v�V)����FJL���QS9���R͗1��0�{�پ`6���J�6�Em���|M��5���V�+RC�J�B<�v`���9dA)�J��)t�~�e_�&Iv�qT'� v�B�������v�G��;X��3������8�|J��d�%��E�R�D/���m|H���G�$�W��#��/s&!�M���!���gh_��3/B3��ַ������w��R�kk"6Fr: 	ԩ�)p����%�u%' `��#�9Y3x!cZ}��V�@��U�CR�P$��՜A�;��5��qdT1�H����rucF/z_����l��t�S��)�]�a���m�����!�ZE�7��sF)�?�6\�i�R�ЙB�����~-�}t%�����2۩�hc|Px�^�s��8�lJ	j(��"���?��{� ��,�!n{���ð؋kWԳ�,��Sr|p�f:�J0��5X������>^
B>y��K����(l_$�3����OqP�Cu`�2��Xz}l��q��������{�����@9b���JU�����^�ڒ�`�,	������brv�SQ���������6��}���>�����i�/�'c����^v��Y��x�ڹi�BY�-(8�E��Ό�(YƇ�����'DC�Bw4 �������'P������*�Ǖ�{���F����p-oh��Q"%���=�:��*����EzlT�,��!n���r|X��i
�O��P��xG���~��߶ǹ�+�v�"VN��o�����v�8��olo��E�D!�P�r�����{�,o�#h���^�t��ޣ�)�Tq�W���h��Ƃ ��c��P�q�o ⧙�kC\�WYŊL�3�L�इ�<FS�1g2%����M;Hy:j����yZ�_ۀ�ޡVF	}u�?�	��z���V���1����#����f��k�6D��(����1-�}6��tB�2,����a���6U��&��o�}~Bż@mP2i�ͩM4�(�QL��y��-�&��gB��"�ML��0�diXeE��V�vJ�ס^�^���h�8�АjX��D�a����Om�k�5�y���7�r����kM�E�O*=�g��F�mI�ְ��~̹(��_�Q�%=�W,�!���@-�o��@�::ȓ*M��J}&�﫭�p�����st$E��J*���M���8�LO}F�ۑأ��Te�d�mh�;�*h����G���g-ͮ�m���r����]̨nڑ��S��ay2Fo�7i����~g��� .ìvVpѫ�N%B