XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
d�gXMR�����ݣu�]�@�5V}{��Ҕ��+�=��@H*!y��v@I�-V�j�cLY��6�]�i�D�c:��4όJt�B���i��Jz�L_���,sg�����q���I^�"o:T���ݐ�:������8�%1X�x��!�%��G�em��J@�34n��a�SB��':�ެ�S� G�����%��:}���uQ_����#R��bw�Hu�1�$_�E<�`I93���g��
��e5�h~���u�r{�'e��a)�^I%Yj���]��?��jCj�	�b.,��h�mQ���{J)��$�biک�L��~#ϩHtJ�1&0�����3�m(�<���]Ai��[��!V^5n2#�Pm��ZQԀ��:Ab�X���i@Fm$�L>��L��*C���בz�~����-+�%���"���ܬ��ˣ]�9J	�}�v��]�q촉��?�c��N���j��KKO�ii�d�ɒ/�u�cK��nG��[qmH9�aҿ���MWQ�_������N��4@+V7VxT����bpB�#'#^|�U8��)B:�����#�����-U�;�gd.��&��fB^��Xʌ���zLE:��>����T�n��>a���&�j�a�Z���
�ط�����I[��L!��xϱ=���oY�쪨�сkN/nͶ�{�B�~(PS����3�i�������ȭ���Rk���u!��V<��|Y@�)Ǿ�c�}U�a���o�mXlxVHYEB    fa00    1f80��(����"���Rw)�3JV�ϩ�g���_p����a?���l��t�ɜ�w�c�	���h4��(}U�O��{ĩ��O�_֚�mOU�A\�=#�E�¸b��=�՚��=@+l�௘0�0��c�x{��%�Mpt�\m8"l.7�4����I��Fl�G�r�q���n<ց�a��9@t�5\���F��1;��G��*�oTM��=#����:��U��n�ڂ��6ܻ�T��_cڈ'c�â��+Ӌ1�=�����:á�&p(0� DZ�:l6{0��Z�'}t���^|��V��C�%��,?���B�IXfP�c�֢����U� ߅z;�կ��oj��^K��W�Ք�����.:��`^u�*SԠZ���"�6bj'���8��
����/��x��4[�W�F�"gW��>(T.�+���
g������fb����}X�����l����>[-���8W�8�)��e�y��<�\I��B�}qe?��&�v�K���ϯ��6�`�NO���:�?�.����f��u~Ho��A7����Ri�Q�I¨��s@s�Ӟm�������rr<���u҇��fw)�p��y<R�E�,imA���$oX@�^��.}�F�V[���6�S!N�A  ��N���;�	q�W���)~E�;O!�7��ڱ:���Z�#�8As)��{Y8n���WA2����:�+��Bsx�M��`�ybG�J3!��ټLZ�O� �Z�PwQ�7�AE�{YSܥ��N���b�f�?��)8wB��+�cH��B�x�{c?�p�*�l�i�Z���x+���*�)��8�&�L�雰�O8�
���Q��UU���u�qd��DnLp����BD�/�X+*DLv ��Z
)�;)mC��u/L� �
�=ۼ��(\���L��a��: ��`i��z_�����TvJ /YD+7hE���8|`q�F����5�Z]m��@�sSY?���Fm�k<YD�L#{v���p���R�����A���l[�|ة\r���?x~e�m���_����?�0Co6p���]�'2(;�H��.Է���B��'�9DN���?#Z>t�����M����en5&W��ʜ!G�?̏�U����V3rI��OT���1TM&)�<����m�S`�]������fϝ�Y�<\����VFt���63\��Ĥ�F���L�'�����G�Z�*7M'�Ս���Uَ%����Z�p�i�#P�zO�&�<V�r�S}G��������ſ�L��Ჟ��Mb���sml�kq"��d�J%qhb"�1��$!��p����V����{�)�~�!N��IU��U��aX��swJ����=(�8�馅�ܾ�I���V
����e�q�r3$��Xb��.�
c��x�`���U���Dd`f٠8�Ҳ�܂h�8GNo�v�j���7M�'	�ԣ~���|z.�S�ɺ����g��5���>�Kz�ocK��	mU�~W��7�(��~��a���p����2�>N��(�^
���V��P%k�/s���[������%_z��O�^�?�Kg8�ü<2H�P�S�h�P�uތrt�?6�s�6��C;�ݸ��#z�&+[W����Ը��W��ka9�;�|Q+NntMex������x�]��N��9L\���?)�����/b��<e	`��<���) �|Z�^E��W�,�tb�;�Q��D`�w�:Q����,�1���Ě��Y��]�?����g�U{��ݑw�rcr �b�8@�zS8�
$i:������>W�#�ڠ�;?�&@��O;x��hM5���e%�@�V9^����ugs����*HG�گ|:��=���&4q~�RAC��'hGk��6�N���b&aᨳC*�	��䆖-q�=S*1�S�u�솂�x�:�X�k��#}(���
��e�h4?��J�P���Ȉ�)V��������>
��z����δ�K��G��<E��.���hi�05	J��5��En�Z�n6H@��G����f��G�4�����_'�Oٜ������U�!���-6&�P�67^�����ۣ]��y?E<�f��LXmZ��.+����ـ�28��c��z��=��_�q��"��J�W��o ����D��+ZQ�R#=����Y���|Sr��a�y�Č�o��B��7���(���Z�%��d��-�SpE��� �`�B%VLm�lB����}ZR%�̐��0b�:�-�ҹ�dJܑ�y����������?�#�HJ�\sH�&=�r �^o�*��*� @�I�!�X��t^��LN����Sb����N�jοc4xmQ��M�*����$�v�^"��n������!kO��ꪤe�w�7���5���J�3�~���
���j	�S��1�S��쥤7�l�EE�sT� �]�y��,�B��s�=�~Ж�9>ٷ��)�z˱D�%u���ԇ� ��m)����t"/k����������7���4Y KA�;�ӝ�����&��V~�!�ll�ٝ�u1t߂��m���/�	�i�yDbkW{^BxN�s�8���dQ��:�bM:� (@D���+�d*S/�p(2EC���� �|��5Y7]Ĥ0O�� >���Ë�q��6r�w�h���ljb?J�T��m�Km�w�d�fE0n�P>�å�NҫH[� <��|��tZp)��Sl���/�Ej��_�V�&��އ��Wh�MS�H�ocB�j
�o�\Rg��rKgwh��Y�*0K�>F�a k��yJ�JS���O!�|:�ލ�	��+�a0R�2C�gF�0����Rz>s��K��X9k�W(��AGe��!Md��I\t0���9��M����3��a.�]�¾�ݚ��A��xc2������Mp���bz
�
Ǎ�@���$���y�&�I�o��.Łu�M8S�����
[~��S�&ǥV��A>�=�Ԗ�wk{�uV�U� /��A��B�������@���9��k��$
g�u�#�]�?�h�O�p/�g���js�؜� `=qܙ)�Q+��^��0�O����zF�0�mE����	�1�F�Cm�A�rf�;u~qPB���s���eW��lZ�]�Zd�\����1Ŭ"�0�q踋����á���Y���AS��np���>��z��p�.�Tfz�N<$��I����=Q[9Z<��4I�7�����{.����3=�u9=��́
�?��]d�.���I���T���%�'�����[����%�}Y_��Hȗ�ދx����7l[@��dGe?�DAP*4��=����y�<#{��v�~��� z_K��6|�U#'�������=���Ն� �g
�I�����RWu�
�L#f�D�9{�W_��iu�޹.I��vY�
�Dn�����FO�1ڹ��G��-�����{���d�b5M�R����}ֶ\�6�_�Ws"��y�@�܆��S):��L�[m&��=�}�#�F�E@��>l�)��Yz��D6CDK �0�.�lNAx+�dR�����������C�2*\�-:`�7b�Kj��	�j}��L�Ë���w��+?#����37	��W
F�խW�{�m�D���[�%�3uV)�Cgђ~�T�$��0M픸��gg�������U�_���~��.3���ǔ���˓Q5ý�w��4l�*�Oe�)G����T��k�A;X�p�I���b1�K�ضj(o��;)#�c�P�(���s\��3V��~~<�Y`!&Y�A�����������FwR�H����G�E��9:)��)��G�$�/�Or������Y�����k18n�ˬ�]��`��iflVP����,���ij��l�EBW�v��N��2�Dץ��dh��W
a�ͷh!���ۍ��(�A凚��u�$(��O�fJP�J!i�Z����w�ZyR�-�w�+��Eƥs+�1��Wg����&�K[�gJH�̕�s�����'�"L�9�Y2��tO�^J\Ծ7�Ǻ�aO���`ӥV"��\FmF��+�5�N५:Z�8�����/"U)���h�#��>ɼtU�0Hx?�\��ռ�b�ѩneV�L�VW ����C�;A�Hw`ԧ����^*�W�M�V�LBg�tt���Y� �{(2T�[�ߜ�V���`�FS���	��M�3D#�A)�"��
�Sa���"�9t��$�z�.�h�^�j�Y���WjY�"]L6;���� �_\�q꘶W�X�H��m�9�Iգ�Hn�v����Q� �`����"{<��'�}o�������~ok�<�	�Vk.��F��x!1[U\"g6�:�}8���� 1���F��f�.AϿde���P�&1�dX��5_��?D��� ���ō��@ajY�9c�n���2<Ƴ�ST>f�'uz�K�j���C,C����e3-K�o��ӗ$[��ڜc&���m5�j�"Jx\�O�#��j�NO�>�!��=��A�n��q>�Y���N?*@�����؉����rz��<�i�dZ���}����{��ۆG&��-_w��c$�WQ�u�s������9���1�fJ%݃�S:=��X\�,%��X�����F97�o��fE�w��i͜"zY;jd²߉}� "��v7�D8�(��\H���k6�TIpQ KMN�[LEN�	_!��rZ�v+-�s����F3%`��]VY��t.����-s�(R��冗�r1.g>Y:��E�����F�wT.��z.%�|��P�[n�L����*��Uп/��tS��n����k{�84-������=����O�p�d��UҀ�	����"N�9l؏d:� c)t�7�I�1����wim��_��~��#$������ �;9>�����{Y���� ��3t�ܲh�_�=m�k�ƴ_��s*�
>��K�Y7Γb�W�5ĕ�?�3��W�n��Ω�jh��Q��j�!0�3
��C��� �N��,���U�Sث��D�<���`�/�K�T땽�j�J��+?(o�/}��2����8�?����p���qtzz�f1��[�LtnA���9�"�}{����C��	�F~O�`=,��}enf��j:�����Uf��U�,ۼ�;[��ay�H�s�'2U�ۧn�)(���b��^[o-[��?ё����T�og��	Ã�W��o.
�pĄa�&�8@n�y^�ljnK1	\���y,3.�~���I�����lc�WPD⯡ं}C��nP`���+QB�g+ռ-ަ�%G�����X�D�vN��ɕ�Y����GO��Q	�m�;��QwܭlZ���p��"	��ٍ��C��7K�uyZ�R�W�h���>��Rb{PUh1xǬ�ܭ��׿����j��+�܈�ܣ�;��2�"�~��y��M�_o��cUϽ��4���L�w�-��3�g*�UE�"n��(����55�{�/���q�(��5�L���}��usys~��w����Gq�c$=������w%���Tt~/y6����O����NFr��� ׏����P�K �1�X^����ئ��Yʣ!jǵ��p��߲_IP��&{V�#���
.j�ʭ���l�����bI��l��FA}Cr<���&�j,3��<w<�K͔��lem�F�q;Up/�6+��
x� 
V��*��oa5�"B�"7,�>��7��?���νE1�(�i���jc�B>~��hl��\0 I��8���hD٬�9�����P �p<v���5���X����ٖ^������x��������^@��z���M��qH����6��6%3O����Q)~@T�I�$f�y�?B�{�fJ؉��h{�=��U�����!��{"�Ĕ�Ø�g�s�1��,�6լ(��Y���e��տ��>:��&ϲ��I���C_+�@O☔XV���.�GS��`��Wp��N\'ژ勵*r�����)�9{�?��ǀ���uఠuo�B��������-��TJ��Q�A�����6b	��D=!w�c�ڝ�T����qx�l��;p��Ej9�
4h�!�Y�g~s6$��TG��6p��n�/=�U�R�Q��m�=�na�n�ql�l��AъPہ��QL������5.��jEthg�qt�BeZҺ�ۨ���K2vB�.˓v���^����Fs;K��V	0��a;�(���V #84��j|p��K��+%�ߖL�����Q&]�)b����Oh]m�X�Wi"��KU� �(U��M~���{�x� c�����ꎷx��\":I���?;��T����+�o�Zݤ)�9c�i���rɧW����!�����v�{��c�[��F)�v����n�)VY��UI���t�k@�[*�;/��^����X��*H��� �����4�k�����Pt+Z����+[�I7�Ή(��@�杌n�³V-�,a3�K��Ɛ׹O"s��~&�]*�:�ܟWr_��Gn [I���6JgA��DE���kMX�׶��_�/>:9�W���6�A<��L���\�ʊw;is����̎�AٗJ�����ʝ53�j�kY,��F��Se���p4���h���Le�҆NV���眱���X�P��!���N3�gK$��v��uA��+�
��b�E�wS�߱=0�����2N���ß֊�oF���ߞ,�v1������ �}�:�c#8��#J��cE�+w
j*Z�w���+�-�h�|q��c� 0W]G���6�!]̬s�,���tq�"g��)V��ʠ����c�����#aa�� ������ߵ&�#0TP���Lƒ����띣�g[�I`���IK ���3.{΂5����qbG�P��خ���7�t�6�o�Z(CfCE�L6���҂�P���(�ul���C�Y��۩����f���ߎ�E��Ir�';�HJK�S������?Ga&�g�o\�EQPJ������GA����t~��^9KāVZ���ݳNۗ.(yH�@������K�z9v�m�%�#RF��=��m�u�����B�o9=Pڇ��?�����1�m*:�+�4�4��/'E����2��<�R�i�&71��}V��=�G�V��U!J���9�<*��ET��}O�6�=��W���<j�8P�� �Bp�`�-�!��H�+��6~ډ�S���������١`���D4]`��I�A]�li*�j}����5��H��^B��e,���λ��g�^ (9R[��>^G| �%Vf�]����m/�z�LΞ�\��/GG�|,�i��,�heA5t�B�];
B���,v�)�j,(�{��'*�
'�����,������]�H��9)=�Rm&Xָ��7e�Uiu4o>{�������OY��|�^v�{P%1�q��:�,���X-��5&�g�2=0P����u�q'��X�J�K�1T��Pgq}��n������m��0��i��e����$a�q�y��S�`U�+��w��+�,=h��BV�,;��p�M��Ț���}���߽x�g��t}Ɓ��C��>�`�!�MH���w�)y� �g��E�BD ��Y��-�_�P\H���a]��[��B�P����itW\u�S����[Xfŷex؇�R� ��[ʧl�v��Z�j	��S�ٴ�aޓ���2&�Ȧ�e�=��������ٽ)FPs&��!���_�,5/J~�������E�~�Ϋu���la� ��2�-਻�yv����������h�����{&)@l���C�2��ȑ�@p��1��#2ۡH��XlxVHYEB    fa00    10c0Ç�;W��W�̈�4ZA���l^��x�'��\�+��pĨ��7��\Ȗ��&)%�e7�������ֺ=I�	� ��BF��j:V@��7�L��nj<��𔕪�v>%%�j[^�=���Y�©�Q�.�
�M���kgV�t���釀R��F�(ԏ��i:t��u�Y� fj,\ln����!@�f�֑�lb�_�_�7ୁ�4ܚ�_
�
��(����#�����������4��牱7�%�8?}]-KN�2;Q1Ռ�������g;]W������|Z�U	/����l���6��<l��ͬʂ�IܞX�r&l�/�0$�ۗ9N�����h�+������
���y���)����������V��1�<w�98�Y�=��=ϱ9� ���P�pJ��t���H�dC��Dp���Q�2XUȉ�?� ���N�ǵ˰����s�qõ|
�|9�m
��C����L��5���'w����E��9�����dUb�z�i���P���*c�w��đ3�ݤ �����zNβ�Z*�`���9F.�^��Hv8�g���fk�ɏ�qj�5�%C�a�G7
�l:����97��S-"�[B����Q�t�2*(� ��`��������O�Ƴ8M�=R��ҷ��M�*(� �y��ȝJ�Ā/����xUԀ~��*0ǿJv$U�j��*[w?@�$H����\�E:	��Q����{��Ew��)O�ݓ}*~(sdn��J����Yр����~~�TIu������D��o���n�g�]�&Z����;�̭�+^�*�L0c�AG9	,Nu�x%�|�3�X+	�' n��	�t��
Ȍ�*6�*��e�$�	켪Afq�"����b�ۈ���깹lN�8��Լ-�E��I���a�@�d<��ùj}֍��xQԼ�P�Jcv�W�I�K����M��0�A�}�
-�-����(�j� ]d��b������s\�
�k5��T�jI	�HͼB��`MJȷr���+#�6��m��"��ae]wh�R��7.5��"�&�\AtE��<�p��K�K,�g|��������1(�o��Hdu@�����������Ô��)ڝ�[|~ju����F*Ϝ����):l��.y��h��w��5nd	�'`��ܕ������A(O>�����*����w䀲.׊�JwЦ+}q@k=����Np�7DG�z�d�&���0�^$#ݝ򡫫�)l�����W�-�!�E���� �8����Z�yg������)}��R�I�y8�%�#J5�x�y�C��jӵ����BZ�,�����'Q�.���S�Z�g�-=0���t*4P|�)���aD�V:�@L�ԋ�Χ���d�2��������(<L�V�4H��A~����	��sng��J�� U��%�6r����B�`��5������'���~;ZV+lOu�\��m��Dy���a{��r��[;�)t��J&WV/�ގ�z�mƇ�� 7�9D���L�P�~�ߐ��2o3���]�����Q��D��i%B����3S��<t�����n�����)4�tJ2]2������W:����\FD]Z��4o�t��9c��Zy�C����~g��Bh��Z.�m��ݤGh�[��F�+��wyAs���2O��ܴ�Iߜ��:ec��W١��~B�T�R樾zߋ�|H�𶕜{&��{��{��2&�A{����9�H~����>P��G.�\���Y�s��O|GC�_C]��t����ʽP���V������+�B?p(�Dٝ���@�p����S	/��9��5�+�#��E����o�%��-9�5]K;�˓���^�!��P����{hT�4�����;%��wO�o���F:0y˹���N�k�m��S�%T��� :t�d"�Z�}�N���ҟJ3�����̂^j�A4��nfp�>��^s]�Қ|w�?��Z��ǯ��>6GY�~�,2��w|Ͱ�~�'ʲWK`�Ȭ%{;�{6��[���z�ꯖ`<w��Iy�BY�c��0��`����[�Ϥ`y��&>�nr�~WA"��X1&АR*���� $e2���'D\?�?|']jAug P��ԫ��V���Tl��,s�/'J�{�����ʽ�I���A@kA�o�X���� �	�����\`w�ڨ���6#d
����IK��0�_=$�S�ؽ�ci�x�w��;`~��� |.�*E�I| :n�Q���,����zu�����p�W{^�ui�3k0gl���e_��3]�"]���<��=k�+������������P� �Q���W���[�U}�)�+���a��Pd���鲜o8����ֶ�������1l�D��j�v���:T�����C{�@�^��V���4 w/��Gĉ�G XaxQI�h�4{!����VFQ�� 88a�Ѳ�"H[��֢�xr���QY(P��?� �`�v[���(���0��I�\\�%k���Ơ�!��
W�ԍ-hrY�����wO�N�=�Gtu�dv�������q�A;����B��t�2�.�jV�MG�BI�ؿ���+�|�2���H��?�K���=t ��VbE=���e �����=��׾�vBޑ���f�6ԛX���<>�9`9$�r­�uT��q"^6�q,�g��I�����:`����Xj^�Uġ��@��њ@�lZ��

� �~	\�g߿u�9�������|�[�����)��7sE���;*�Fօ��;;���l~�ؓ08�"���>&[�Qc}C"m$�6!H���uy��ŭ���;i͐)2g$�Uɘ��<?�1��VG���X�u�o�'�Y��EhU�&H?�ڎo�32T���O�_҇T��|�� ����+���Ω Y�~6`����r���G�T�.Ԉ���?�-�q~tG�u_�Y_W9��zY3;��1SYr�é�H�=1��ӗX���k�vV�����k�Z�4�⌯��*�F��?[���wR�4����m4�ި�{s�tr-�O/1�u�#��CJݛo�пm:�Y�X�W��΍f�� Aen����w�����팇�L���0�k�^4�}P�px�`cƌ��8�
�_:U�K��y�f�?3��tc�;)�9��n��a=*Π*9&��4�H?osV�������w����?M����q��[�ٶ�
�|Xt��"�V��
���Q7��ѡ
~A�
�/��eI�j�QD\�ڥhm��3�%�|��S,;vc�E��&[��쁆%�c{�P��^*O����I��p2�������HP�>lG�L�Q���G��翥�����>�#��k}~�B���l/%:Ϊ���w�K7q��\�R70b����$0_P��,7���7�$W-}��R<(u��S]�dv��e:�ݯ�E�����7޴��R��1��6kw�p(x7#Dr6""�j���9����wqQ��)��.D²�w`��q��R"8�}��Eg�y��.-q��K�m�t��n�O�HdzcB��t6�S5	�X��qu����E���6��ޯ]����]�����E�Ȓ���� xC3��v���j��$�Z�_��}ڽ �M]�/���P�@�������΅FSS���7�nU��/<�P(��J 咆Q���O��{P��(ܣ���t�
�������\u:\�w���ȼho��8�k/0u�/���w�u�1x`%��_%d \cD��Z$��n��+��=D-/|���K���Y�����Z�'a�T>��f��
GW.����]���t��t��ͯ�k�R�dV���o�غ��O�W~��^�i�[�~��#�f:(�(a/����C��Q�)lkg�VզXC�暻�Z&-�'�6޶�nz1u{�;�k���\�h3��!z�;
�ڙ�͞�1�u���&U���b��`U*�6�Z���h���TLo�vx"��G	X�u��[��n<��k�����ϻ��Af�a�jD�W*8~�������߱F�Lh�~�/k=�,�{�8���y�x9-�����J��ycYgH�Kѵ&y�j"ߢ�����m�aW�6H�-xf�P�����ד�lH�~���ˎu��AYG����v���͈��rE�e����M�)�P�'7<�L�P��S��Q	�;����@��{�#�tU�����&D{5b�	��-��XlxVHYEB    fa00    11409�.��mx����+{�[df�)=I۸��3��R���f���9pq+K�R��*k��
��oM�+�:�q��4�N.��F��AײH I���������mk���#��t;_�^��.>3��nx�r�E��S�������D��c��Uf�D�q$���蛅��NU:�ۼ���G��$I1"���P���Y����ufg�!{p�P̙���i���4�u.�h[��H�"o�����Z�y7��_���º׾�W �<	����J�!�&��$n�x�/�[٩MA�*£�i�������(j��1�0��*���5+6}g�+.�ǂ�4��/߭g �xrK�
�%8��-��z��'\~�U�w/�(��v͍�_Nn���fDiQv%��Ἇq:���8��0�x� ���i�o�"�ŕ�!����bhv}��Z���������y ����@�:�`R.z���*߈�@I~�1@�*�wg�]��Ùn�C,�چ���3�&�WfiO���r�=	h�D^�c���ք���\�̪k�a�����A%N��C�@!��C%#�M�
�}*�S��-�+��5d������S�Z��w�:'a[Uƍ���\o�^x痳,���&n�n��#�l���v��U ê����i��aو��ԉv�j[ǰS�>;g�1��N�|�ID�*d�2�Ձ�
�����sCvӡ:|����()���O�b7�4��ʹ��a�<&2����<{�S�K��8�vlNo	.�K�\��4d��ǁ��z�F��M�u�L����lυ��_��:W(Q�Fbsʙl�(#ak4 �!(�D�f<=�}�S�cߡ;{�6_%��qa������H�.�s���~S�mok���l�8n�3��k	u���S�Aߖ3����X6��@�!5��<��|�O�iEo�����l_��qR�y��nD�sIMN�k`���\H6����X�xҽ�p2�=cN��[Gר��H-��O�g:���RZ�ٸ&�9��멗ݽ[���I8s��l�Spg8&��:�D ��<\,L1�sW}צK��jv�,%a�w�(���4/o4�Pg�^�-����W�B���'�ip�\�LH�~���MRh�䗎��S���u�3��/~<��l0��Ce-1`�=SH�i�IjО���,�V5�.RcÆڒj�je��!1|�E���'t,�@�"�e���v�Dٿ��7olf��|>e���@;xc;�eV�F��y|���S��fnpͪ|c�*����O%�c��h���b�ю�ރy��	 ���Ŕ؉ڦ�=������=��A�q`�K�2:�0��T��B�X/������2�QEJ_���r$
NA�9 ��!{B$�%Ԙޙd���Tvr!{I�u��A6e�&��PHͪ�v�Kɸ���t�7�����J�6>� 1V���0���X�Z���l�]�۹�zK��Cz��֙z�m�0�6�1s�ٱ��u��R?D�s�n�O�=BmV���?���+e\�Y��l������U�[�T��4ݥ����w������᫧�����`���oѕ70�<�'(	ё�ԪS*I*=����'�r<�NJD�_���,�ۃUٳ�IZ`Gj�M�B�~�9M�_㭍�}?j�R�T�׊g�_��^��(�)��?�Ά�>D�7�@�}�x�<���U<�:��*���˒o�qg;"�J������/X��[9�� �^�$�+�(	��?FÁk�	��R9���>{�t����gS�6�ٰX/MP�ĦM� �Y�#�R���_D���x���8�n4�B�)z�b]�D���<���^��-HN�r�ʎV_��҉��:�w%4{F���(���������p��_d�E�e�gA������-S��=z�����i���b�IX�F��vD�x��6B/	j��u�fQ��˧�O5�����EVЦ����A���9�$1������C���_y�
.F��K����Ҿ���W�bUdY.�����a~d^�)7���Kȕ*���+�jI����bK��s@-tΐ�>��#�}+�L��Q傫N��FP}[�@SS2�B��Agy��4�\���Q?���Q��c��s�yu^=����� fV}[j`�!�������H�lPŬ)NV��qx�W%�S��m�q��L9Wp��9�]A�S�J��[	�������$I�12���F�o�R�G��.��J����������ͨxk'{J���حK+@Ӈ��Z$Íh�l� ��W�j��dz�i�/��hktL	׸�^�Z+���D��t���k�a�q
��-;9N�0+�7�v�Ⲹ!6E�zCG��y�!@D\N��c�Z���D�9�k���Z�x.d��� eY���u"�cN��9`����/$2��#�ۧ�d��@L&Y������pJ���TQ�n� �\sl��P@Z�-ԫ��P*�{�W�W�V�˂Μ�G�pIS������m��}ۏ�/qNu��:v��V�N���
{����^zP)�~�8~�UYCxΕ��4�ƵuQ<�yZ^Di2�3�wk���p���XLp�$�c�4K?�L�\c� $߸e�ο��{�7���6ط��y��0c���G]��V�1&e煞.��Xl�ɮ���t���?�K��V�������3Iдw����'�z��]b�}��ʟ�WV9d�k{k#�؂�	��C[��f��{�M��&�8 ��w�{��Vy v�D N�yB��*���,�|�Y'A���R��m���>C��(�V�N�����ˇ���"��N�1��:Q�Ύ=�QY��˵O}���Gw7=��8�&!lc��1"��@[
��'<�]9޾��W_ۊg�D)(�!���s���11Z��&ha�6�Yvr��ˇ�Jk�h�P�K8�x��$�2�i*�8�k�P�oζf��鈺�::�`~��qJ<��	��F���{Z�A']5,;��[�QT�|
�y| ���&������w���� 2�̓a�:0��V��5��Pnɧm�����H������so������e_�)��G�����2![�dG�ʣ��);iv}�M�/a�7�bi0ۿhRR���7a�_���LUWM��Ϛ7H61�4lh��
,�ͭf�ZG��i.	r�Zқ�&+Ӯ$���]�ښ����?���A����l���2V��/Z�H�dde.ԑNHFyUh�w�cz���}{q/g�5�p�X���w9�2��0�h�&˦�@�0A=2�)a'�@��Y�S@��%ǣ�7R6�&*�P�I4Y	�W|6���3���I��ݪ��č8���B?Z0��Kow�;@V��%����9d��h��= 2}��G�ָ"49���_�u���d��+o�#���y?��)�!jT�8��f�ZW��W^����:A�%���D(N�N�
߲rv�HmjE�ƙL]	32��}-� �hԐ��HH�h|�2Ũ����У�z�����>b�ޔ��;�����j���
���Ď�F����0l�$(l�asQ���.��H��¿\�C>���R��Ȑ�5�o�x�MO�[�N�^��Q.0��Nn@��`VsS�
�$�C[CnĀ�����@�r��߿��r����f�/�#S�$.�o�����fL�>! ��l��%�3%G��1�(���M1��y�_9�L�U�i�tr�w�1g�1���)�kݓMl1�7�٧��a\��*�����vh/�?̥`��x����Q�#YV-��<�9�mO�Ҍ��6���E�`�N0Pª���չ#��Ⱦ�?zs�`� p%�1<m>(n/�x�5��+�_�j
�#&�(h�æ��;ML�,� ��>�#?�I��h�T)��L�r�M�L�&i;�?���tv�_(��u��â_���ϣF���OڧA���"��䦵O���E��b//�Zo>����)�:V�������14\���on�})�dK�Cm��?�-�=�psz�&�9��3�F�6�Z��X�}�Y_��Y�e�,��?R�u�3���o�v���^��FW2tU}�mBTl�^b���������̙T�ҀY2?�D���xm<��ǖ$�[/KԞ:�0�m?1��)��J��HvHy�r�M�w��u�'6p�'���V?(U)`�RSd����G�"j� ��'������n�h�Q�^�4C�toɉ
�j��������$�Ꙣ�$������=91=���%�:+�����(>�M=,T�=�j�����0����T��&���h����t�X'(���I��������6�qјA<P˳q��;5
3��a�XlxVHYEB    fa00    12e0y�����E�X�Hj�����u�B�)�x8�56�zJ� �	��qfƋ�u`��,�2����h��V[߹��(���J�}h5��A`G�Hl�Չ�٧�����x��J ����a��nӔl�AB��	-]K1�z��� �����sRH;I��!9��~�R���V)�1�]��r`��Y\�=��
����9��?G�1An3��o%Uk���gq���&�FW����[����I,�yˡxvp�L��Q6��M��6��̎�*��F��1�tZE�s������F3
�*aaE	4飏%3�+���ƛ,�	�ksr�8ҳ�"�b�)l63<w��S�a�Uw�xF1�x4AP%����JG3��{܊`��C�Ǜ������BM���袜��ؠT���~��/�����֟�張1��O�h���DS�No�ŋ=;1�J1�)�t:'�2�8�U�l��~%����m7+b�i��F�,5
�����FPR�	O�jě�Mf�����Lδ9��/}SA=�S��(a�YqԼ �^u�fИ�k��Z���$�L��!	8�v~�J��q�43z'�r�o�v�Q�?��P���;;�`n�g"ф�.�>A9C������u^��1Z+R1I�'HR0H�)�����@gJ'���w��B����q�&���@�9b~o˂�v�Uq�.�0[\�זJ����x6%�d����K�e�hI;��t%�f�
4�l�(�Qo��N��� �Ƈ�R�mE����eb��5��|U��	�Η:h�q!?���t�-�.��$b�L�S��"/궦�ܮ�n��v����=�w?x��g!�i9���S hn8ë��Xw����bt�؀�;n�G�r��0���ő�<b̄�R9nŦ���s'ًD�e����hu�T��~�@�'��w�ک-�B��lD�r���� T��3��8d.��f��ԩ嵎�3Kh��מ�zw'Q�X�/Ts���m���{5a��WO/v׍���a^��6�-��H<>�.��n$Ju*7	�>R�p<�yo���z�͝��C�4��ٓ��Ұ;���#��PP�����@9�Pt�s���uƼ;4)�L���� ��SC�u	d������IG���.�'�K� �9 P�|�Ҭ��:xw?oS�g���_ժ2A!�[>�D��II�g��2Y��7]��IN����SԢJW�~#��!>�+��b;ć xm攪�(�~䵛�vP�v�9T��C�5���rOt�W��O���_�K�]���7�F	��P�#���UpE���+;l������� jl��G�t/�%Y(�Xw��x�R,}�A t��;B:�m�ȴ�[QEe��LH�+����3��&�ࡊ�׎�j�bA�T�2@����Y�r&�嶒������T`2�Ȍ^/U�����;xJ���f&`]!�*�U4��U*��.�ᝐ��;��i�S^ Yx�P��H<��ƺ�R����o/�0�.��E%���{ߒ��p�T�!�E�#~��JXd{��l��*��zD�x��M{Eh�
��#F�'��(nJ$�͆ֈu#aZP��8Y@QیFFމhh4�� �b����#-V#7ً;�C�^�7�����b�'|W*z^	!�2zt	��v�uS �s��%#�<�>bb�)R�iG���I�����1M�������˓�	疣{�<{��z~�D�˨9���pFǅ�C�5���3	b�8�����+�{g�s�/�DU�?�ʹ*���=/�n��q�ۃxw�q�U�+�ӟ��`��������u�R��j�%���������A���Ơ�sԲ��3���_�!�2�����2�Kө%�7>�	�1�3�׆ɩ�a��[��w�������v1{��5T��8!������|�m���e5 ]0X�s��(���/���:J�
�a}Ɉ�B`�+��&�����g�xw��z���Q)��#>�<q`�����}PWg��v�O�ޗ��-���M3#�@l�E�Q�����*Qh�Y}���鱗�Y6C��q��,k��7�|Oل�b�������T<_Σ�?�����=���wW���������x�%���[�),����.s�R��4�-�.�j���\æt^�)������{�3�$;���b��4�&PY���фkOEz�\Jr�G��h�;G��ə��:@I2�I݉�,@���!���IK�:�jE��wਕY�x�Z�׼��yP�0�JIqc%��w���i��h�\TM���a��Ɵ��}�Yz`�wQK���v�/7�>6�+�+X�;:%^L/ʍW���jX<�M���E�3�6�G���Ԣ��$Q>��G��ŧ�4�J	z����
$Ig�>�*�/���� B-�ݴ#:U���G�YW�G��7D��h6:�a�{��P�f��I�T��e+>��V��Bg?��c��Rt26��tT�W # �8��Vs^�T����yY��+��m�b_孱I�c��/��zD�n����*2�;E��߫Q �Z���@��tS�ܩ��Ago`Ñ0	��<5�H�ְ�� �/C�B�G�a���s^��q�/^x���#�K�P]�{^�;(-fj����Y_
y�|
��!���[�����G��J��=�p�P�xڰ�bGp]��1�UW�f�yEh�h�7^0�:,�a7�̒�W�S��-��h�g���A?�7��h$w�
���ciR��(���t�6MU˷w$g�}NVPǌ�;��7��|����d�;��?]$(H4����E���U0�Xh�_8zB�
ɧ���3U�*jo�w˔L|/��8XV`��Z`��;VVV�&�����Y0"��`�Fz�#�Dq_,2K��j�@�7s�� ֱ�=L@aW��MSzGKӃ	���F�I�2�$`ק��	�9�Ʒ�n��X�h`n���v��ɫ���O�� .�$���E�:��C]�ڮ(l�L���{	�N���>IdOx�)p��A@.��u��*pb��&����,*�:��i����.�s�l"Ь���#<�����G�O���	Ȕ#�9og;#i��w�Ry��}�z�r�";������5�c)�&:�9vܱ��k,�Uτǥb%��P0:m�*S���ҝ.rN���<�&b�~ :H���
�ô��͎T��|d�!���t��ّ��#����W��-h����q�G�n5��K�H�nų�A �6��Y>h ٱ�Ծ���^2��T��4拹�u�_�-览} r���Aq�oxGa�Z�m~� x�A��� �Q$~	�b�w�Yŧv���lM;�
�]c�!o����	V␌����>=��S��H+ku����V5�U�	|���Y�j/�t[-�B�xN6�E �qV�N�w��4u�������h������������ݻ��.��<�.?����Rr!�<��ᡡ�D�z��=�ԇ��g�xl1J q�ԥ��m�V2�����$N��a1�E���� '޿���{���>/�][�8��7�O��W��My;�Ȑ���b�';�� �R��T��Exh�h��Ҕ�Y�[}�V0�gU���t���Y�F?F�@V��5����Y�_��V�h_D]s$i�]a�>}Y�yl���9P�J{?߰�����,��%��R�ڙ|f��f��ËI��I쒩��Ψx�8��a�0�V�CT
C����5�Iiz�ˌ!a�5R�yo
���펉�u�࿗�v�e�G�R�!| �W>��)Vr�T��J�/u��ŹC捉6O���绕�XN��)fэ���UL�����k��s�5�����=���Q��Y���M{E�ٳ���8���B�HIm)�G�^�$,�pi,.c�m��!Vd���:j."���� ��UJ�(�xz9�>��"M	��J���!i��(����e�R5t�G������\`MP����s�&�G���`�+���3��Ƀ���ת�ȸ(*���`jƸD�lI';�D���91ϖ�^�w���D��e�����}'�RA��/f�͋������`%d���k�2��.��3KC�gaRT��ۮ�V�C�f��fc-�M^H���y������F�ds�z�9����_�A��CJ��Z�z0��"���ͭdv@"���;Wy�x�����#���hWG�/�*��C ۫?ҁ"�,�V�Z��4����J�]���A�r�@G/��?s ��oy�/<jo����9�'�d���H�oo@�Ò����^�Meʐ'���g'A8��|��#"��O��q��T�?�IXk����qM��V'��_���#c�=�����;��B�}ݜv7=���lc��޾�Z������+���?E}R9�*j?WӟDQ�w���O�zk#�Ȇ~�v�*z�����?�����4��9৴����X�}�U�P���	��O�+��3���JL�E��0�yQu'zccd_��Vb�ƞWuwθ�}�lË����|ݮ��4�ֹ�`�)=�+��ʁ 5���K����V-�8��[\'v+d0��L��N���(M?�F��ԅ9�޳䧖O9¼�����m���A$�l���aA\�Q�H��M�ă���UO�?q�~h���vG��98�쵀�����FH3��	���/�����lB�<�p~��M2Thw��Z ;�hfXlxVHYEB    fa00     f50�T�z��=7�Z��R��Ѓ�*�����A�4�a|�s�ʑ[�E5JR/�嵍���"?��!��V'4Y_d?ej����t#�J��e�q��q��R�<��.��m����}1��O��i��!�=���	OAO>yЫE=K����b8�RIn�As�[OC��ڨ�?�<���Ŷ��ɠk�_W��=[C����K���-�{I��V�c)ly�m���jy�zÚf3(�#
~طVŖX
G�/xena7�o�'#M�V��΀�U�δ(��y����z��%t�#=�Lu�
޻�̽�����(�޲lr4�Ô`�_�ʂ.���g�����U��cS�	x���1DlV�dvމf"j�瑀���[$ZQ���;��Dy�
��0�,	0�7���;,+����z�D2��b��1�a�7��s��+�_�|�2!��]	�>va�pk�E��N��,��.�Y2]XD�tO?�i��ؼ�������Q��	�����f���ܝ�7�S�Lf�1[�a�I�_AE�D*ل�6���!�d�[JN�'�ĩ�Bq.�bݨK�T��4	 �M�����VJ*�Bd��
�<�J�E�3w#v4&��I�U��9�í�2#b�Ts�T^ �g7֮�R�����t�μKc�f����<`����'����������zJ��)K2ԟFQ8QK¤�okO�w����p��l;��t����JK�}E	'��Yp�iJ��[��`4)eM����z ��5C/��h�"+�L�A�񄁁#hC��*w���>�_x�,�X4�@����8r=t�/DL��3D����<���3�W����<o5���o�m��L�r0��8����q�^^��|�����R���P��.���� �"�YӾ/?(t �"�njiy۴a�����:��I-�7'!�1a�*|��7�˫o�z�������{�2�T)�:�Oh��A���CX����0g��A�ĥ7P߉�cA&��ȿ�O�Li*E�@J��X~|QH�d;����b�`��-К��F�Z�����˰�
��螯U`�.mMANCx��h�OKs�?�E��7T���j<�tWd¹=��n���ɠ_sJ:�$)�&�����o� �a���3�Bi��^>��uV���&B�2�3Z~I�=���_��菮�*;+�[L�z��q3��cwt�rn�A��i�?�b@\�x���P}�R$�v
^<b�v-��o��d@�v���g9%�!�Pܮ�y��.�9�ނ�G
)�>�.��.|�:5n1vRy�+6uz�R�؏ 4��v��a�<z7J��{���CJ:�1߽�d�%���ּ���k�u�S}�����vYR}�ט����WT �Y> w��g�H�f���Y�@rH�
)7��4����-����.4�@�C���Ġ�5	,i��=u��4Vlħ�!n6�,��.�c2}�>c�}�Q�A�g岗�b��G��+GH��b@$�,;�x�-)��~�`���&#�0� ~���Fi5�I�D�hrʯ�8M�� +Л����*�3�~���y;�,I�8K�(P0ƹ���f�^�n9ڥ��V���:�y�k�N@�UOG�&�Q�c�D�
�SE��-�o�+]��孿j:��y�>y#��N}ϥ�JQ%��w�:�9O�{h� ����?��C.����ɡ�}�I�X씧��kW����;[V����v�jI��~ӭ��4��6Ĥ����I��d�x�W����/��
 a��+�����3������9Xhi4d��>����4Զ��W38�����<YC���:D��4��k{�c���t�F�+t�+kH�+��tRq��u��1ʌ�|hH�Fo]�A�J@d��J�c��v��󷚙����Y���L��Y*�܂a�#o75�dh����Ə&�KX1/Ɉ��Փ�n����6�k9����, �<j��� լ��T��kGǸn&y�=<���t�ډ(�i��1���i�|��>w��?�cM�/3��5+j�#�͹K���'�]%�:�f|�{�^�ݤ���p_����BjB�Υߙq"'j�0�������vjM1�4(OW�ڍq̴,�*��s��`���ϓ�6�Oz��u$z���0���ʆ�
�@m@"|I6�j��
��;FCpP�6xx2$�F=��V��"���a�N
5��<���Sc��_P�Z�D-%����;�Q�J�n/��U����&%3CAe��dҕ�^��N��:H��4�P���2�C9Z�#8匾��gV{w`��.U�����\������T���o+kH?�[�~��A=��7{X�@�,xfρJeb ���^S^mQ��H���X����r�����t���Kx�$�\, +?� A<�}���wi �`��_�|���Φ�[]�kwߝ�g�q�Q����\�F
�?_��`�P��y7�R�/5�f�����Χ�lW���Uf���|�N��9�C�Kס���(��-���xچh^����_r8�OUI����L�4{.�Pvv�<J�{��D�X,�\�Qʬ�f�Z�׵��R�+����˗h%�_rM�@��l�ŀ��с��S}�7W���?`�I��a�9r�Fe3E�c�g��.0�k���fuGG����7v�*�&R�����k�Ah7�����6%(�>&ְ~�i4���v���c�����>:�||h����*)`��N����yUɬu
��br"cLӄ+�<]i'��'��o4��(^ ���܏Q-��.�	2#���Ӄ�=��s6��	��t��h��*�yqqq��]u��'Y��_���;Ԫ��.�CJB���"JϠoLJ)�;�QD*[��?�����lj&�,�,�-��f��
_�����"�7)�ۊ�iׁ+IA���RV�C!�u����*cR���I�Q�R���S�Ywr�W�h�[VdŹ�~�y���j��k� �x��I2DE! ���+O�k��U$_�z�=����SH}z��� ��Tj�H׉d6���$���YP�g�1��^��1��w�N���\���*��*BO㱆֓�K�A9�����xaӞ�����
i�N�PV��;��n=i�cB�?D�5w&	w4)�a���	3�Ĩע�+�u�
�4x�W�^�ŅB}���w��`�����񓙋�b���z+F��0jk��k�ǩ�"Jo�r�j��O����sD��#ha���,FO?ݕ;lQ0�G�/�	��
̏��7z�.�m[����R���޿�����m�r{h7?Z�8������o��|ԝwc�$H'���n��V�,D�D=�b�H��1��McqS��[���L���+����7j��W��`g�_�V����+�R��7�8��}�ȑ|�~�K_�_���-R��F�2%ć%	���E��b@ݔ����u,�>f+%z,��Mݲ{ɞ������>����[��pz y������[�X���8X\���!���]�r�gpP��5%���b&����zMT�f˭X[�7�'�U�a�]��/I�4��q�����Ms�ox�n�%&S_��� �K@
xE�P��<@�߱�h"7>U\���aH=���s?�&9_>���D[�1܆���a����<�iw��SƼ@��Nۑ[7�O�{K�iwE��{ļz���OWkB
z@2
��u�0�>d#�9c@=�B̴�t4��Wh��4�H�$�j��<��o�&|�#+}���r�"����:�7��������L#|�;�Z<���C獅�������Z�R��^�~tFT�1fr=���g�b�ǩ�VG��&�A$�F���p�^�XlxVHYEB    7273     560tL�<���*/�l��Y�N�|`;���P/�_�,%����x��x��by�_``,SB1��"�G�����:ލ�r�mS�Y�(`筻����	dQ�V}:�+1�LR�xD7��v�W�;=�����}-��V��!,7}I���?���Q�GT�f���|܆JS{P f���� )Ou�+%J={���:S�0S?��*&w]H�i:��P�Y�ƞ{�ō��M�5�G�B ;w�k��ښ�h2	y4ߎ=�13��Xecc��Bݐ�P-�w�(B^�ؐ*A���Y`]h�������$
e\���_��G�Z]��O�6�fc� ���u��z��r̼�\�''z�Iw_��5F� -�/��W���1��o
�<���]�����\��D3փ?��x&L� F�W:+E�Q3#�#�9�$��7Dm�Ы�j[5��(#�	-k�������tD�Э{���~�<S����b�1�0f�aR
c��k+�]� i14	,?��-aO{Q��.�w�Aݑ/u�������OӘ�FU1�pp�D�W���5eM�������yZo�G�2��+L.� Х�U�0s�T.C̼�0Qz�Z���V����i���i����N�nH 1̖f��e�7���`t׭�8k�M��D�5vtwB4(@꼓>�o������[m��;\y|p(��r��C��N����ӑ�Y.>��\�;�VY��+k����k^���b�!#���f~�Q�ܗ���'1Y��c�L��4�W��겎��8;�.;�|�j^�KT���^H�#ժ�vx��ۅ��M%̀V>֡ys��΁�l8�k�1����b�l�� C')�]��u���)�8@�t L�\~�_�<_�O���2c(q:_Y���1��p߅�����ڕ^|m�HV�p`�;a���:���`�1&��sW�辆�_g��]
��pS�`��Kڄ6GUy�A�9���U��/�ѩ�鮜�9@�$��y\
��<���t���?��<(Yg�f	�۠�+1��wC��J�JX���,.qK"�gE)e|?:�m�dhD�����tZ
Ҵ_�AB�e_��!N���	~��9}�8�8�B}n��뭳P撝����O���$L'2���+��v���S�����h,����y�����)��8d`�Z�l�&!���(`X�2��D9+�PkmI��ם�[H/
(/���2M~=����G�	�6�0̓`���D_�X#]i�����q�К ��3��N�c��<SKUS"˗y�4��JK.	�>�EݙtlK�'/>f�y�2�_����$ƭ�l�Մ�*D*ʦ04�Ax*J��8n��#R?h�S�*v֭