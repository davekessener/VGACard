XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����30YM ��re�%k�P����x��Ţ�m#Va�	5��Y�-���:>� �39;�I�|9���
�G���YҒ�����l�����m��_ҁ��5y:�SivBM8�B�Yfv��=�}=�v,�?�;߼�_QV�-�5����4��޻�]�k����$I�ȍ��m�e��D�9I�x���jͥJ�]N0�b�PZ�v:`G^`�0�T	O,e�	� �O�M��i�v�M|�7 w�r���t��q��@�#�I^'���=�LEcgF��gj[�J�,��F.�i<�	��D/�f���xF���Յ�E��ގ�v�� L}� dn�ºw�u:���v��>�(�k�/D��
�N�}T�D�k�e8��P���E\��ހ=;:g�B�%�8K��Z�\�7dN�i��#�����~��kG�b��3zVpX���jI?�Zh��p�-� J���0����}H��Y����W��c��6u1u~1P��N1A�A����|��}���Q��v�m���S����W�M�L��#����r�BS��'��ŉ�*����k��<:a�g'�p�a�ka|QNV#q;֧7)�/�A9�����B�Sx�/u3��ԳwvS9����[~�K�e���'�<�Rr��ٳ<�R����6aw��y@�P�B0�9��$��T5��N�N}�I���j���<S�co����9��[�Cq�D���_3���H4&<gͭ$��rvX`�,��&�؎�ݾ	$��l�>�XlxVHYEB    fa00    1790mU�w��&�t�"�D�H@:���IH��-@|�-�ڨGƠ�~�T�D?`n,�	t��ٶ���,�Gp� [��K`bU�h�^ٳͨ�}�M����놜�����V�c4Õ����˓�2wy�m��$�.�ط
����ed:�Q��R��A>���ڀ��`1?��_�D�L����{y�-��Ѯ>Cd���χ����x���Y|�'5W�<�]˴-���}y
O�M�B��MS��f�G��������_d����BbF.���$�㙪��uJrƿ\N��ث�w4�k��GS����h\E�R����ZQ�g�=]�d1�����<�;�DJ5$�c� �1���D��{ T��G�P��A�ƻ��hq�D�C���@�~Y�G���u����_!����"��b��m:9U|���7����~b��Д8�a��F��:��u���$��lRT��`\�s&a�������-`��p�T�8�T�vō��e��v,���K��a����Gx9��8������{� ��+{� �a��A��Zt���X���c�.�h�tprxe!P�sX(�&l2[|%���/�$ރR�UB�e�P<P��˨/���7�j['\���g.���կ4Q��75�ʬ�<�r�l(�gB���7���*�����fy��"���2׍M�_S@�+`T���I��zs^���VB]���A�j����Ӵ'�$x�H;���FR���}��W��`�hx��-,��r��
DÑ�,������/�a��/
��l�_�sH���tE[|��k�N�{���H!6�䂯�C{�}�{��/a�I�(���晟0��h_$ɽ�]�	���=���^�2_�6�T�?Y�8�t����@:X_�X��V�;�B�IŇ�Y�/�̼կ���[���f8̛/�\�����} +�����~Y�p��w�ZI�7�!�ʙ�IԊg뤱(��tdcxN����L���qS^Çx�C�1����D/�`�F�m��$v,T-�4�0�Zm4`�ޫ�<�zڂǃ���>G�f�jRt�����e)��\�>�)*�!�H��>�SV�s87����"'Y���u�7w`i_,X4�
p�}�_FJ�mK��)�����l�u`�W�@P�e@�v���w"�a�L$6�� ��v�I���@�j���^P9�m�U�_�?pPc�>���Ȥ{��K����w����\O�S\ղ6r����@�..��n+F��f��Ռ���`�7Lùj�{��R`����+��@�\�_������2\����a�gg��M�~��R��ܒ��y�B㣑��E>ϊ�U:��"���&��p��Iˋ�Ø��]�V�3�r���RN0��Y@��7�����XzG�	�>I���ϸ*��-�A
���LT��=������AD<FWWd���7���x�տZՒ����Qj�8{���o��!�o��=V�M�ϧ�kyH:�ĜH�5��ъ���5sG0����}]�2�/�0��T[�c�/MM0�1p�5�(Z�]�,��Pլ:Q��[ �������J�r�@�����zF��`�,��ya��u��a�aON�����J�De,��cAxy�IЩ�%S�k4H��Kp�;��jC�M�{�^ߢ����"l��xc��:kYo��G{��-�l��:��57F�� ����E���(���̃�PQ�OZ�_#���N,������}ba�LΘ��׬�)_�(��m��%���݃?�WS�n�r�x靁pG�*������v-SƯ��`>��w�;�&��;IϚ�����]���GF�)j��T����_Nh�u[)��� :`� ּ�C���/>�i�ul:!�.�crO�r�͌�Y�w����q���+N�=�G��M�p��7��cpS���7I�g����*~0�.�y�n�y�:#�*��&J`�H�����������Ֆ\�lxHԻ��׊��ߛF݋\�E0/a)�ԴLZ�ٞ��z�i9��]��ޕ��z+W�f�3@e�׈�&ƀ:|�+�{l��e�z���p<U�_FCߚ��g
�n%�zg]Ki
����;L\bհ��E�@`ƙ@���o�[�e<����\�,�J�O
����YJ��jS�ʕ=��܎V�0�RG���+	f��B�޳����"��x��iA�F�@�u� �~g[�ib�����u쀪uu�W ��M���51*eL���Hdr�\Q�sbX�5�}��C�Ƣ$�l쪵DvJ�ɣ�=�i����.�ǟ��RLW�Àx�>� �u���Z2⫭s����yU�����3�.�C���ҙ�X�bɦ�LV�]��Oɥ�Ga��1&T��l�������獭<�YfVhى3#�J���gY�}�N������n��p-�5�]�I�d��3kB*Z�zM �2	��´�*7z-$��a���E��d�r��T>��O������ҕ������5[ي�{�u��瓞����HI��ѽ3�o��cq��܄	�r���=]:SO�c*�5a��زr(�]2��!	f��Δn�U6�N�X$	Q�)��i�<k�\h�=���,!C���r"ɾ�O�eyK3�ʀ�s+HM,{��#�e������k$����gnh�Z�[~�Z��멝��^[o���r�|V[���W���L'�B���W���/��2����e����!$z!I���q���YR��0���������'�_3�JW� /lbو�Z��{�V�,�(#(x��H�D�7�|�!���R|E�[�w�ꊨ.�7*�Z�O>��M�pu����s[C.�	Ĩ0Q62�b��w��i�S6t�!����E ٞu��je��[�6�o �P7�k��?�7G��
v�H�3�,��IN�(��i�S��w���j�g�7������i.`�p&.�R���8��@oM�"�����kW`E��ބ�P��o$����`� ɪd�/�D��O���0�y(_[�6���4)��Q��iM��U���܌\ E�yJ� ����3F�\�G�vY�:�NWTU6ʽ�(�m��-���-L�L���T��6U :����4c�ޅ��Pzfh�=�B�$�D#߆Ö�)��9��{R��D$Cu&�{��s�^pI���#ܩ�V�}B���5G�B���yv����A?u�����V5�#@��/�ϖ�������g�m�O�ئ_��:��"�Ph��b0����*l*Ǣ��EU���G��u&�Ϗ~7} �2�v1��c��۲x��	5:����'Mjħ<HeD��:/��7ގ�Y'���@�%'�����uQ]�il���2��MtSq4@UI�U�������#o����q���vF������	s�����4-�v��]�I2�X�5��"ӊ�CŔ���w����8�G��Wc�����$4ܖ�H��bMv\zՌ&�Z�Ә({"�		罯H��?�U�d��i�Z���r��0�Jk]Tt�3ȶt�\b#|U!������Ծ����Aخ(DGb"�B�M�L^��!]>���	�,�}:3{	������y$w�FF`����r�b}�8�;�ΪcXK���!��o�P{���c���4��2���7�98�ٺ��FŘ�L��|���Tb1Bi�p�q]�<@5�ΐc^�� ����_�S7ݩ�jmk�1�e�`��Cg�0����ˎ�؆�!�����(x�$�i�&�CE�'��x�h5�}U��@z�?߃������ϱ�I�Pl3wXH4Ҋ�"��(W����t'4��Z~�EU��j�h�x]O]0B�Bjd\2T٢M��u�.���	s^a2�����89v2J�]���8�Y�.��wRK����AΙR�0d��
��lf;����;������w�r &}�{���k]`�3�A=�o�$<Є��:U�7P2w��$�1+l {���&ps5�	�)��G��a���`��f����dQhK�C 7��:������OiH���@d����=PoݠA�9�lԎ�)yZJMmx��Q-���iGH%\c��-l���CQ)��\���1�"���l����hA=�:I$�N$4��^�Q8_)����PV�ӳ"O�'n�4֐�a�6�촗�w����?@����O~0n��=Ћ�&ŷ�M��$`��BU׺�k��5�~�J�y�W7o�o�ѺvֵW�-m>��*wE%Cc��a�y2����<��칣E�g�5N����jO��h��xv�L�82�Sq�����萸�XIgb&�s>��x/��~��������i�G ��M����-��y䛒ƇE�%��Y �τG�-޴}c� 
��L���i�=o���*K�L��d?[�E_s?�o����Ct�1�x�%W�Y�S��$��ȇ�|�BC	�a|^.�uw��=2����n®̖��zd=�B�5��|��[���- zv]�.�j��77v���L��M��V�B~��B�%8�4=��&��r^z�zɰ��H7 ɍ@YJ?��ن��_$�Sl]��+3/P�ߴ�hD�s�ȱc��Ub
2{���=�v��LDBGv��\��[N��u�JL�����b:#c�M9n�G������O�N������!��m=���p��82�I��x_ƪ���U@?r�3��Q?�7�R~���)7�t�D���m�$���u�=�*DO v�z�z�>=��p�"������
�a� �>X�<�Cv�&ũG��w�M�����iL�Øh��1$Y���Y��T���p�_�wX���|�	c���Ef`�n�"������	e�G�����0�����c<�6M���v�����:/L+'�f/����+�(��ѠN�/�[�P�����lg�CY%��V>̮+���-�$������l�B��;vΤ��>���]��8b�5<T���mĀv��[�3�%ϝ�Cc=��y���]�s��
RW&�#�`���g@G���S/=�(H�I�w��Ro�n�L�{��t�c�Rҥߧ��8�v^��|[/�Yo��%�H�[����p�v�=;'�l47w6�JB4�! �[^N�k�4Mn�+�+?s[/]��z6�)�-����X�+L����^Ȣ�Y9�����cF?����t
�W��F57�z��r��@� :m�`D��-$����!z�G��`6���d� b�z�@�.c&���ApFE�ɜ\�h1��t���sԃo`h�$~St[�S+x/��o̮�&W㬛-Ӛ�똄��l�ex�z��j�M�);!�i�^�Q����Լ.��T�a�����n�ø8Hq�9��`x�9�w^]�{��A�����Ĕ�AUQ���؃Ñ�'����4Wꪙ֏���V��}MwGl���g��Ҳߋ`�A���
 ������5�a�8�f�
���j�ΰ{1wi����qWC����%�G:Ly�.�=��%V^���r9)s�(�K)�I��0=�U�|��{�C���v�mG4���k����	D�H2�x��zZ���{q'�H���B�=��Kߧ��5Q���� �Ȓ֤h8�YI�1�c'&��|��}䙆�Εz&W�."x?)p/�e*�2����yI+F�D~Ma�}�q6��$����2f�
�" �ns��:7p_��[�f[M4�ģ��f�Ne��>�3۲Vg��R������/�Jڶ���T��KQ ?Į)��F�'��1�X���]3\��D��&�$��Ш베Q����Ȥ�OD���a*�ΰ�:���y�?�>�&ZEn)���>6������(6��a��n\)�������i�jf�Ѓ�[5����B9z�O��@T�����D������6C5ϼ����f�G�#k��Z����/it�����w��kF�[ǘ�K�'HXlxVHYEB    fa00     5d0����*&�`�:��� s��?g񕰬���Ԝ^�������g�w��W�t�g"����~�I[-�r�%򱓁a8���58<�JI6�p`��E@m��5�Fq���DGvG5h����6Z�@IX��X�!��wK5n�1iO�>CD�V���:*^H6�c��K�E��ٗO+%M[fE�ܜ�����q�4/�ADN�J��վ���_�'�fV~��WEs���T
���տ��5
.�vȥD��_��*�z��rSL/P3|4z��(�#�*�wW��r��aN�0;MOI߅51���� T�R�b�����,џt�JA���^�=� o[k��k��a[ƪ"Bc17�vt�����k���6�1覠���ɨ�}ޞ�]{�jѴ�h��!hXʐ�q~ٕ"���:1����͢�PU�YT��rm�I6��*<�n:���@$�X�L7�]u�D�.��9�W�.I�(	��2���q𷏄[Q�X�I�g=9����� �
��D�t��5��(��z}������.y��m�cA��,��ΔT��?����I̳�]�O�1�"�s7��e�^��o�����[�T��"�ҝ}f���=(���+�cؘ����=���%dw�<^T�#�v״V��6!qx�SN,{���3|�]��ֲ@�����U����؝�ڼwt�vYl�&X=�3��.�΄���.��R3��&�6.��"���a8�!��+#��d:xތw'�~��Z�Pv=2�4�8^1|4/x9�&̟�?~�$��˚���O�vۖ���'H�@�G)�u\e㌆�$U2�ׁ�W��8D�7�[k��t`���)�OA*�E7���[��~�uؒ
��ra��9��_O'���:�M��m�����-�'L��] �K_&��U����8����W'��̢\��Q�D|:u���q��ll�d;2�T��T1s�ڑ����b��צ�>L?']&-��<���S"�	*���֌索
+���+xc΁AX�X����N�'�H��v�k�eb�F]7�����(MV��㔗����O{�O�+��}�Ä��h��O�N(~n��)��?]�'\�ok�*�d�� �]B�
��s����櫶��S���wA���S��V� ��B��|/Y��:�;�-.ڧ@�i�D(̩���|����Jm�^8�b��=5i�����u���9���K`bd�2a�K+bl5��/
]&=� ӿ}]�Y���c%���b�����-V��� ���T��o�k\ʏ�%%O-h���uۑ��uU����.�/Lͅh[0�����9  �< �:� �j�S?9b�<�Fۼ4طFj&"��-��q��o�IPrx�J�cw�Kc)�1i�_;}O�M����ڹ�?�!�b�T�c����;�AIj�a���GGZ���y���=��8Θ*�5�r���X�XlxVHYEB    fa00     640gN��:$Թ�����S�7b���i0�1&�	s�����\�s3{��&6Z��8U��� ��-���$ė�9��1�5s�����:y�k��R���7d�;,J4��;�>7x����mϱ�H��P���I�P>�{@�t{vCZG�X�.�.h8���Ү�2Y_��.2<�ۓ��]�U̴������H�b�� R����{0�1���4�,�f��	�5�(�X%��=�v�؄]�/W�΀#]�G�s�{�!��@ţЂ�7,2���R�=z�.���(	�ca����&ջ�VG[�_N_@�pA;�'p�:+^H��a���������.W(L�E0�U9}s�������g�H���e�9�5M����,(���pW�:�J��I��t�+��e#�c�yE>�l��W?��j���G2`����l��0EF��w����A��� �+4{H4�O�D�u��	j{]�aƧ1/�%��uo����6�UC�n1�N&s ��[`M��?
�ɡ��1I,�(�E>b	��-߿�g�y!DM�2�Q��zb�=�ok5Χ/^5�s��6�n��ߜe�L�����m��S�f>�|�"��w�-VKG��S4��m[ܷ��+���"8���r�/8P��j����:�w��^�a���ݜ{�+��wa�'O�|g��J�ڦ������u�"[�'�Ӑ�������c�d�O����Ͷ�,�l"��Y���t21TW�Q��r���1b�A��J���z��O�0�������Q���0�Y':�}`_�����ݵ���T�E�a�k�����'�m���{ ���Ҙ��)b�̳�� ��H���P2�3�PԺ܉�@3�d�Bl@Ȟ�"=%.��N!'�zN��z��k��i�~*y	�ߝFͳ�'�c&�D�2��W�KU����Ad빞�(���+ћ��0jD� ��L����WǸ�t�n,�56����Za%�<Z�?[U>p��Z<"ZuEw�v�(��V��@���h)E���lP�b��ϩ��Հ��W8p���/���qN-�g�.)�f���u�LF:�(Q��;܍D\�WR� _G�(f6����:�I�@��H���tJo�t���v.�S0r��=�_�aw�<�� h�v)
9���(��8����z�&`�`o�.]uF���)�w}�K��@���R*vo�i3�(V&�?E�����Ǚy��R(Wp��)���!����܁v3!SGee�c�"��B�������8��i���}�T&�m��9fS]v*�����������Os�����~�w�q����j ������� O�ޞ�]ͪ�{c��[O3I�F����*(@ΐ��N5.�[}����X�����Uƀ�lL�2НPJ��N80.��dw4O
�<+f�ӣ ��p� �-;@�(]�y�l!+��xs�0P5��/��j�+Y w���Yw��9��_Y<��!���9vc���L�����q�G��ON��Km���N]���z�*w�ҽK��z͘x��.��M��Ț��K�X���jz]aW��;���<L?� �k��XlxVHYEB    fa00     5c0X�M��ff��5y0��ig��GU�������JL�й�Ǭ�ipv"�:�a@}<�v��{�[�.6��,�=��q�a��J�[��xS�!<S��ďk�B�_K���Pe�`��"���2��$����X��3�=S0x^��{�a{��"	��K;Wf�ie���ϜB�+<�] ����5;�'�t�G�[�@d�����l���E�D���S�N�_�Z
��	A'��꘧*x��ם-\v�$cW�)3�..�������\�����4�OdCǕ�m�L�i�H<^�Ȕ�a4\d��s��ׇ��E�a��h�^f3�/��c�n��t����Y��~�x�*W�Sf5�Q� 1���1�4C���vI`�+zV{˯���#"����@3�-V�1rb��uDo���KJj:���ٹdepQ6HZ�^`�M�������5���%�8[\�kN[�Km}3b�]s�~܎kV�&�~��[��U\>~�@ˑ�?i��Ĥ�� :Ep������C����o"��z2�]��ʜ�.�=�
GӃtq9ih�c-����<��aԽ���Ie�5�Ž��h�x���or��yĉЏ]�k�d?�J����w��|��y��F�r����e�B̵�$�"X�`�����F��g�d��u���Ŋ��ɡ��`�0�9�rҶ��f��f@ćBRD�X�?;��M�u������Y�̜?"�g��l�i����g~	�;���b?�HW�I�@���A~�<V�����Zz�3x�H�~��F�(^t�:��4�x��)>_W�aS��:�d�Eآ���t�S����R��1�Rq�ʑz�1�S<,?����\r��|�S�1/D����/��eR��XψTE�fUT���^�U�Fh�L�L�*�����E����$c��܇����B����c�1��߅H(��/���LKL*=���\S��(`ˊF��NKZ�V��>Ub���=o���0ؿ�Y㬁��GQ� L�֯�7��A����C��G	Ӗo�u|��"E�����d��4�xV`�r�к�݆��:p�͖of�E��-m-Jg�eHZ�{�)��d�>���]����t�D���3�D>%n�g�?��US�Jbw��"x��`�X���~��̰'������u�f>(T��ۖ��D�w/u+����o���!xz��c��[�HM�C��P�A�<= ���)4�2���nE؂l�W��Y��1��ڤʐ�P6�K�+�@�R�`� �X��HZm��^�
9�⇝/��3gK�Q�M�%nn��������5�iz���G�xY7{{�a{����xE����`0W���?pUl;)��E���%c���X��8�8��
�L�fhg>)?fmZ`g�r�?a�:`ᝉ�D�kp�Oyj
_Q�-Z�:hP����hC@|*>�)9{[�W��:=[�XlxVHYEB    d347     a90�C��O�P�ܕ	�g*)���7#d�O��RcD�j�i��]�&92ta�>�	^J]�/R�\�*���ܺ^��g#35� 0�Q'�T�8�a�l�����=�7�H�\O���z��T5ΨU<�C�F	��S���4j�{�qw߼�}��x|�a�R@�B���Ev�藩���m�أ�] �Po'[eiǳt[�~�CuSfg�N�%U�ʊ�-�{����N� *�i��l�cC*�� *H78����z�u�>�����xS��g��F*e��W�YK���[X�=�O�g�]v��J�9n<+".�>l����i�"x�������F}Jj���YU��	�@�)[�*Yx?���� ���G9�at~K|xw2�*���F�^ ��?)�c6�WqaF�q˪�8��ʌ(f����7K��Qn� ��hi{���f-/�Tbb"�e�-`�>��U�����I�\�F^���K̈*�P5���S*-җ�K�02���I�|�N�PD��"T473Pѩ�=`��3L��ђj�����n�.I\ӅFE4��\���M����l�4�-K"�[w+����>D�����_.��ݽ�&I>Sn��])�Yj�ގs�r"�t�i+TA��V*T�}zE��޻��;t��N$�.�rc|Dx��@���������ͩ~��[7iI����/��r��־۳�`�-�#��V��R[�&)���D���h�sB$�tk"h�)(c�fx_�_������.�t��o��]tx������?Aۗ3�,���=�w��Y.U��ר���!�pFHR}�Ox���s�n�qtܢM�� ��F=�h�{6�)�'� ��@>��<u�C��H<��%@�ºUF�]m������r��-`���(�>>V���2F�p��<i�{�0бZeލ�yޢ��;��Z�]Vr+/q��n�i܀���4vK޿@�W�g��]:��j��Xgd�2�s��륒�I����Sb�8o�f<�Y�D���t��.Fc����њ~��G�e}1�\��L]&4RU<���XI��
]�,�����d�.rN��/�'b|H
�:64c�?�(�q��g���3�g۟�ؠ�-�.lq�C����i1'Be�,�zu��/؟�m[�s�$�2����p��$�S`r�	��|�0"�y���D�Ӂ���)F��M��"�}�V]��B��η[L#�������Qh�1c�{Y)ccm
r=#|�����y����:�/��#3_�0�@���'�'���?;e'o�㸚��%�`��E� 6ﻫK�O�Z��_F�L@�{���xy�,�]y��L넨�zJ|?��O�zwԽ��e{���[xvJ�a1=��8J�E�ҹ��C�âfR��L��:�Є��U3Y�"�l\,��9�L��PZ��aH���%d8f�@��y�D���� hv�+�7Y�ڏ.�"�|l���N�7�`����ʃ筡�����F��P��Cl}͇VCG�������M�_��1��o}��6�+	��J_�ŀN8�VS��K:����_^a3Rߔ�U����`�$�����c����:�z���L���]	��,@-\�x��;��=����_��VW���S�Oh�NsfjbpJ�l"�ޢ�|�`â�C�D��Sf}NÀ=Jԓ��W��F��,�H`�����a��mg�1���$I��#r��b��Øو`
��u8������n\�q�Y��j��lˈ�_�r�
���,9���	�Ά����|���KK"��ñƞ�k���=O��2���H9�|�@��#��R�{	�ܥ/H�L�����Sl5�dL$��?����F�q.{�&��ɮy�c^z��b�t
ނMB��Fw	�R�\r�j�oHgY]�gl���Ϩp�ɞ��J⻉���#n=9Iu�ܾ"��r��ջZ������0F�wa��Ke^K���&��N���E��\��r�q����gT��/χC�f�a�,��v���w�v�#���s�ю���|p(�7���r�A64-�u�S�;����"/�`o�!�X�I@���ѓ^+�r蔈7�Ȍ��g۶���t��÷xY�ұqKB#0\��e��Q�g��<�f��1�f"��c��),������H1�#�Q5�2��?�
D���	@%Z�F�VGd��+�=��`5q$A�a��*Q=zT��=w�9۫����n���x����i]n|3s�לu����<z)��LU��^`�gv��56�k�]_�>c'���h��
8�}!�1:�f��Y�/-��6
�����CC�b�����4 Q��{벝ˍ0�����eN%BE���rs�[���Zs3�Iʆ����"���-�[9���$h�3��� ��wXy*�p��&1 ¿���v|�fT�-���+ �rSRU#��ӓ�"������)���O���$=���u){���u��HK��Nz�i0�ݼ��FT�x)�:[�>c#����aȝKo]���������
�sQC-��)�Xc?�8X���-��u�T�������R9��k���3�M���G�Ni�Y<n3XI��fh~�@&�e����čܩ`�k�yJ���F\��|9�[���Pe����<`3������p�%�Թ*9��#�߲��~�J=��h�P��~