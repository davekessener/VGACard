XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���C@^�pb�¡�9K� ������4�1Z��}�\��"��=\�A��\�|W@�F�T'%[��W.�?��Ķ��g/�{ P4P�l��pkv"<a�xAT�Cu����΂�O��-=�^����h�Jt3�k���kn�x�=S�	F�򝩠�<O�p.�1��)X�7早j[�qP&���0f����������+�E�1�g�y� ��ZcР�v��*6?��ut���.�M��!ր.�[bZ<���y��-����om�g<p��؟t1!�2T�����v���?xW ^Ⱦ�A&C١��R#j��+0˘lfn^�%������&��B��]~�	Y�-f0(��>ք��l n����b��d��Q���s�(iZ���OS�t���[c V��T66Ǯ���T:_���7Ru�Q���#u�)Z ���H��5C��4�]�{P�o��. /�38�˳�f�u݂��(��.;����tO�c�3V��P�v�=�3�!F�c��8���*Z��5U0KC�w�\�qZ/�k����e�5�J�N����"����%���=��� ��0�K��pW���$d���V��`�f��o�	S��k�+4����X���`g����=�7+��/M�n"�z:�Ę<'0}S2�1�;#�y-[�M�ov�K��y�.���L��E�6O�]R2#w1�_XKZ*�ݪ�a����p@_0����^���؍~J���8#x߹%y�z�1�>XlxVHYEB    fa00    2030b4�0����lģ�MԼF�Xt/Ʊ��:�8p��jг���)�n�p��o?{� ��9�S�������eG�{2�� ��p���TI�R���{,aA�������y��/&�5<��U��H��p�����w⡠Ϻ���Tߵb���Z� oE�>;F0C����/#p뒶��#�"��{����#c����+�b�_�ދ������7'�x;A�etDL�k��rh�{�<��m��v�P
[��L�3���y�Ut:����G Ww��n�F�iM��W�2�B��"���X?$������Ȟ�`W<[��j8�n�9Kͣ׏��_��K��R�?�Ҋp��� �q�!���vߠW�7�ʝ.8;����,5c-����T�ѻ5���u�+�i�W��$��y=c��m�w�W��,�B�����C��26W�����NE�<������Gx�����|_&¨���pN�����F��m��9ѳ�~��[�x�:��`�̕�^������=xrWk6^��αy �6���w=SZZX�,�'x�W:�63t���K���a"�%����1��C�; {���i���٪��)��u^�� ���	�q��Q��C��Lt��A�y<(�9��6i=�E����]��jA
�x��
�K$jc��g�l`�C�팻�&���Z��Ÿƃ�J�漾����N_�9�2D��9I�r���*�5|k��k�O�֤���'�7~��ׂ �2��hQ3�'�)�C��]u�\�\�.M���ޮC���D\z*�N�V���6�8��KU��P�a�{+����s�+uކ�;���0�
�g�B?�K�	>r��h�M`��~1�C��~�R�������}�Ԝ��Q�3���6;��������b��'�D��Q��R�u�f.� ��N�q�D�>3��X����u3BS�F�����Z�Â�(�hK���b��ۈ���C�p�G�Z�zQ�?�,r�# �v`��E���᥸۠�����?P�gl:���m=��v�O����B������S���@����fj���
��'�W��ő;t� ��_��̤�ui6,����^%�Qܐ�N|�jI��uM�������˟�a.�#!2�|N�����\S$c��X��%�o�}LD2C�~b���J7�YPKb�?D&+��+
VI�b��`����YOYd+F�MӃof~��Ԉ��`'#*m9�(�a�X`�N7�'/���c����ғuG����R�����=?P3Ǥ����I{z�XԢ&��� &�� $w~[N�,�3���%UT��4��f�e�F���$�r �����>,e��rI�dk���Ka�x���-x`d���N���\+���#!9Ȭ*sT#]\o޳T�6��^�u���7��D%�1W�U �L��h����Y��%���/�#"o>�~����V2w��zM>@�<|����w*�%'QgL�sd��;�7���1Ir!G�W�)�:�����~?��z�P���تsG$�h�h���$*���q�OQ�pW/zS�Ov1
�(Qf�sm8�m�#"��E����l!�.��m���Wޘ�m�y|��m�(��ja�kv_l{t�����rOD'���Jj���W��	Y�Tݎ{�:��M�	Y�"={e���I[�^p0̼e���$�)�O�hs��R��8լ���R�q�d�)1��#ik���S�~����tPg�I�r�Mү�+�bz�88��i���Y����bJ��m�a��{�ti�Ob������;C�f� �����}�?2;������=mV���@�xC�fK|��;�������*��+����z��-�{�G%������@��j������Ob�P�z=���KU�8}$�E1sT�U!���f�$�t��wVC� _��mY��a����J79B'6���`W�c1�Q8��x�����W�"O���z#�Bf{�K�������#p	���n������@江���e,������ wrop���*0��'�j��&��YO�vhu�&B��pu��0nH�d�f��[�I�/�D;�ly��E<�C:l6�W=�zQ��C�] B����k�\��o�����(X�κ�:�#��������Q�=\k�K����W�|�(g�+5�j"�n��M�񎄜zSI�#Y��J�Ѣ�8�.qt���&,��pm-�ɵI�h��a�S����y��W�FR3�����P�N 5�ʖ �ydt�k*���d�x!d�v����ca
�˨�q�WS%��w��D�X	L�q��fO���;'[��>����:C?�CT�ڦ�lύ��[޲ޗ����,�M�e�j�n�y�~IQz����#��I����Q"ν�b��</9p��T�eȯ�u�3�/��Ɖ���3Gkĸ6>���x�,�V$F�,�{�\\�9��2%w�u$m[m��=�M먖�r�'��������U��}�nc�
�r��4q����a�W�u��ʹ8��'Le����ڋ���b�CB��4k��ŝ!�r�A�����Ja�B�2�B�~; �)f"j��q�u��	ee#V��[��D�g��yK��)C@�m� ����I�-3<�1�l��m5�f<��2��׌J����]^w{�",f�ؑ1/�]�d�7�D���n���M"�T��?)h$J�C�E� ��J���Ə��������^�[jdbps�74A��V��ݧJ7�d�C���D@�aE��*��e)�#n���mS�Q�z�������]�3^w��b���^�5r�C��B!d��!1酞_�����dV�U�g>���K�s�p����-:{��a-���i��p��T=���ā��_Õ&��:�?1�EJN�*9�� 	������d��������[I�M�� ?�E����q��J&�B�\����߮�U�+U*��j+�;ĂG)��|�3Y"���Qx�^6/k ɒgu���Q&���=�E'�����)�r���8��i�X����U�W}睛LM�g�~
����\P�wz-����:�aX���:N�����h+O���y)��b�c�d@v�T��H��f��ƐÆw��kG�s�>Ws�n%������X���D0*�H��TOz�q
��l:����E�@�UP�p��P9cǁ������g5wH�D���(����ٟw2h� ��C¦m��I��^�(�O+
�G��F�0w��SvX>����G�&L��'1z�C��F=�>�aEZK�٬1t2�p��%t2@2{����,%�ˇ~"���	8�8^�u؈X�-9����I=�f�b@Y�A�:�K'��-'_�����f����QaQ �tFn��i�U���o�#�=�]l�`�v���WɁg��n�.�HG{م��}�U��Q��3�-�����\���kKV{����L��(�/Ye<U��dm���f6��,Cсh��2~FB�K����JG�i,�2&������Ua�1�������/z�N��B�iv�2I2?db*玨��6�W�,+	�js�9�z���DL�[�����	�K�՟+L{7j:��m���boMH
�$&p9s�9��+�����	v$�
K��D���$��K2; �<!Q��-�Hjt��FIyX�~��r�G3%¾�n�=�:�O�$u~Х ��1�T?����I˜6!��l8�EÛ�=m�zL�Pj���s�x@'[���QO�͡&�R��</6�ef\oq�R2$6:�"�N�������X@�L�yV�-?��ے��|=-ɦ�:v5�֧,��
*��w��K��������8*�H���WG�@��,���C�U���5�����Ms�����K�v�遐�[:>]�}�gݭ���V,�����˳�y̏�{x�
Gɟm�jzz���.���BJ�B ҇U�Y>��I�_ ��h�D�9G�3��5�u�9z�(�H��)�23��PN�ȏ�5+1�q�fD�E*�*e��?�$J[�;
F�XDE$Sq���==���"�j�F4wNlZ�emC��m�u^,j��S��E�\q��k���M���#	W���*���n�oc�ES0�`~�~�H���s����@e )��'BU�mޘ��D��@D��23�i��ـ7��V��sޓ���+��&�418��3R��Ib�%�����)ӭ)�E��y���L�C����s����!�\~�W7ZѮ>NGk.�£�7�ZN~B�g��t��!�:������ZQ�rySL�x�@�+��ڻ�� ����B�`��U��3�ۻb4���&f[��M���-�ΰ?��*���"�����ѿsN�̚c�iS:�v,�U./�_��j���,m��PK}�������w)��:�X�}�ZS��o%�s�E�M�8�F�'��26�>>b�o�{x�Zi��e����eA�]|���Y�vQ4���t?��M���n�
�ü��ߊ�A�������{��@�����9�yщ�	��I�(��$�=$tYWr��UF�����cW�*�%�X�$Q�6�^a�f��b�Ҡ��lC��i�z���WJcp�'�:�H���Y�H�����^�Q����"w�if��tE���L�>I�)���Vt�^��J�����ͪ�PA�_�̔3F���Zn�6Mg�\�G8�J>m-�6O�K�徫)�C�)���b8$]�Z@��q�z`�nD���Ӳ�e^6a��WR��7m��U���X�1��b��6�ҬQ���*8-К]�j��ֱ�0A��U�ceU«�)����[���v�~����K�8�o��3ڄQ�` �|:zԋ`F�&`O�i��F[�k�d�5�}a
����a!��#q��s֌���o)�Q]�&aqߗٍ�񐕢�Г�ϰ�)��C�8�,�3�ӟh�_��V�2�د���2r��a!x�۽Y�� �a1{ƗK�t�>"���vyw?:*Nz2d�zE�o���6�?oI( 	�n�
XL'aѨ�/s�l�L�%���q�?m�2CR9㻠�9I�R�w�#�/9PLW1��+��PQ�F�v:�`Ef�	j�@G�����8:������_�C���##�������F[~��	R���/��l�֒��Y9~�|�~J��Ƶ���W�kr	q{�8�V�9�� pHȠ����x���l�+��\D͟ɇDQ�Na��0��%Y�լ��k��ݽ�{j�~�A{P-��]Q��4.cX�z�1�<(���`�A�^�|a�Ɍz��'O���~q޸���F{���ug��9��0��~�<Z#��u���XCLV�b�X��=8?�X���b��6�"��U��x���w!�lJ&ӟ��;�#�y�ydk����G�B6�~�)�� ��Ò���F�-���U��ڲ-�һ�4jf���Ŀ��D�U[��񱣋�����j��U�0�v�2�����ܲ���꧂�i��Q��<j���&�İ ]��qH��Y@�IT�-Cث�n#���7��\Jx��bK��g��>"����>Hq�塺�:��.�J��j��E"������[�Wk���	Z�S8���҂�VxR��1�q�>C;IL���8)�8�AD'�'!�I�����	$.�l�V����9��\�Rw͠ā&ĩ���2'Ͳ I��v2,v���]��G��p���*�<қ���E��fĮ��_M��uZ�6q��a��Ģ ��Sb����/i^d��tk@�����gN14����)�Џ���O� �}���X'�i
	W@�ɲ��Vb-��U�G~�T����7Bʈ[y���"�gQ������)�����v'�1'-+-1nN�AО��A�Wr ���a�I��5:�y�YG������⾒��9 ɸ��s$�$Ǻ4�Q�R���FE������%�E��$��\i��ԁ�`7���FA�1�Jƿ���͞4q��*�&�mH�毬� �Z���>���@��엵"$7�n��m��L��/����P[�l3��\�X��;��c/F�?G�B�`2�$T!]L\��h�$����W���Ò���h}�;���1 r�餙7��R���]$Z�Lِ�Z�ڕk�W(�k/�m'��`��3�h(��߯���GCN�lk6���Â��Ώ�ݭ��c(qn� k��Q��D�|���N���9�p*����-L�Wc�7���$��P�(�s��􇫽Q�jO�U��i���jmC ҙ�t�a	����	M��<ѧ#��9s1�ƪ_��r���8��uFF)rC=S2��]�z���/���O(��C��~�+���9�B���-KZ�
�0��x�pn�&��p'�V�4P���f6o�j��YŊ%�^W�k]���^�?
�����~$#����
�u�;+�8�5���
l!p��U%f�~�,;�8���V�BH�s=1�1�%K����w����W�V�����us2��yz�h������O�>&rߌ;���]�`0ӎ��,:�X�b�VP��3t�R�j/�es�9j���iy7x�����m�ԗ�ĭgy�[o(�7a`����K��R��8K����;M�dm6�jSx�y\����tI|�"�^�ˢ ~�`ӌ�qE{x���+dj/���Ic8\:�N\�e-]�B(9N(�	�Ck�	-ؖ��:Ѫ0@u�V�D�m���!<;�A�����
��%gU�i�h�hpC����/x��Π���{~U���`���x���� �S4�i�e��8�8��:�e�����'�!�	�wI�n��;�� a!3ּ	�|)��+-5���Zb$�5�A�e�6\~.�SHp�-��@����0������+${��4$�*�4�Z�>zR�8
��	5��yf��́��Qg�܅ `�w��g�
�/�x��Oڕl����k�N?�W��Z&�䡳3���G�@!x�pp�9���R.~��~D[y�(��罺xh������#� �_FF��&��E]zB��H�k��Y���E6*����C>�(x@�Y9m��gY�ySZRضǃ����J�t�?���v	�BĿ���ꨞK����p�uM0ZD�ؔ��u�����qm�d|Sש���)LM�Ȉ�_�
���kv��b1�o������eM=As��ǵ����8�U9N�9�	]y��r��zĒ�*a����E��U�J��t�b?#x����Yr�|n\�^���*���m�$IU�^����hkg��9z���8w��J^����l����8��>�~����N�|z�穷��2��(�t�T/ԕ~�ń\�%�$i��>�鐁�5�'� X]V�FQw�=�����@C��Ɖ��;$���A۔���m�f�8c=���E�����Qh,W�����PAHŉ�1����nN���G����ti�Hꍘ>h'c ~E�@�8�S<���2��enf�0S!���З)Lm؄��������e<�5G�x�v�f���@��??ϩ�S��E��H�KTf.?D!��u��D�W����?h���V�A�u��g����
�!�gҀD!R>Y�]�uP����:�h��P�����>� g�Л��eSV�,��,	ޔj(@C[ÁY�E�^�nq���Y�3=ppB�f��JB��[j��!��[�+��J�i�(W��Se>xēQ���q��;��a���B�AУ��&և�5��-"�w�w��"���I���߃��%1#;gz-g��9��� :��+��	�~��-z+d�ت�H�D: -y�?b:'EĒ�Y�������F�e֌6uaUy��.��6}^�w�F
J�~�zŇ�����^%�.D]����U(��qo��?��A�ݽH�oC����- $o�1z j��0%	xW��z�"��)�k�9�8�(F�)�♰�saM:p+ʸ�M��ĕ\u�6R��z��v��Q�=�!��e^¨�e��HY��_��*�dέx��H!rF��6�&��ڕ��>f��n����ɽN-��ָt�dd�a�К�{3���2�kԪ��V�[��)&�XlxVHYEB    9620     d70���v�/֜�� lB����5ժ��ˁ��e� %;���{i-���Ap@����΂��'f����sq���y�����~ם\*zO�3t����Ř���>�p����R&P�ȫa-T���F�!y��.Ò��ɥG�����B�"9�MC<�Ǒ�C��>8�@+��+Hv��\�r`[jԭ��W96q�x�d�&��P�D�F���@i�A��D
������a �gHH�3Ͷ�Q>e��W/+�$�T���x���e(�&��L��%�Qwb�|�����A�
%@M���v��Q叜����<�ѿ,����S)���z��|7j�������"S�,zEy:�����9s�xG:�[]ɌIs)[f�\p�7��3�8��co7�;9���ym`n��d
g$J�R6@y���W->���z� ,����0�	�T����o�F�\q����^Z���;�On����BpMQg�{�Po�L�)����G�\X�Y��Ty�ݟݨ*d-�d2��}$�K�u������'>�=��tkEc08���{ ���Ļ��z#�ݥP+uh��}}Ar��:.!� ���W�_tᇚ��+��E9�$"�5xç�vx0�uQ�P�����@�~���ض�s��Op�PAo��$�)����j��9���@V���HrdD��[C~��Tg�|��3[���6����e�\CE�i� h*��ش�wj'��l/j�&q=����q�V�{� �J�Wť�v�2�[��'o�0þ���7ҡ�D9M��<��oy'!n�UNO��Z�d�\Lpƀ���pxq0Y	m�7�LKN9�̉��z~���Zaa�������k[=,��~	������"7���u���c+�߃|&F[٢����4�t�.�z�:U��j�8�d��Z���׉�D��'��W�/��τ���������)e��L��(���ɬ^{����|`0�)X�y8_�&�W�am� �Ie���U]'�fՄ�O�#�|��A�V��y@��
���(��ժ��AG��,L8:3�;���s��)��� &i��D���@	�:�qMZ
ggo�N���/-fh?����ntwL3����0������[����
u'�����F���k�u��8�Ц�h\�޾�NXc�<�류~����=����3�5��Y�M��Ybf�-���2���P��D �;���t�&�B~����H0��2v�����	�b��vYхH_A�ιK#Ak�����b��h����BQu�cha~!��g���F�h}bI�\�ɵĶ�cä��b[i��7����Mǀ7�.����[���5�R�a0� ߧS��؞}�~��5�� C@����dG�_����U�v�R���o�h=1XDh�ʪ`;gl���0m�*m2K@���o?��T��K�)~����~���{��Q�X���R�Jٌu��pRD�vi�{D�
'���#�󉐁���)Zƾ�I��������Q���<MQj#i�:4����� �"�}�֝s8�_��/
E�� �� ���?I�4t������A3���%hI�_i�֛���  kaY�G&��b*%}�Qc=i~vn���*�J���b���� �z}�ђ~�Q�v�MoFU|�0}��M�UW�湻��,��� գ�S�_���ݥ��c0
���*���]y�`�x�n�A��j�mUp��pk��}�ҳ�C]�)�ݙb"~�G�V�>�0���W���x���
�dB�DNVLu^����re"R"hWUZ���,+�3(�d�/��ˊ� ��B#Ǯq��DD���*����D� �[gn�[�ѷ?�&@Fe���Bi���0�#!�r�"�F�b��"�<91��Æ������Y�e�"�	��`�=���o���K����p�L�L�YY&SZ������"X�8�H<�Q�be�y9�W���ɏ���hf��&�z�dI]��w|h�?f��	��MaK�H[B�p�=����C�
G2G�mI�̖��1U�.�jY�3�|����^󂰙�SM��cs��L�0�C��,��u�P����G�����ђ�H��Z�,*��mŵ�v?Ӆ�Ŵ�*�s�:^�jZ�\CB(*���i�6����?r/�EܣW�C�I�Q��c3�ǔ՚>0����2�������G�&>����|â��G�K,��Qs��rVjEφ�:�=�N./S#���:{�^�a�B�S��2�So�=.��M�\�����cy
T��t¢R��ގU�:���B���n�D�	K�w��3l��^l��y? �_r��?�|MI�Ĺ`���P���.L�-~ͫ b=bҦ�>_,' K�\�M�6
l+ܢ�b_�D%P|<�Gk�˂�6�C/��z$�m`���3`F/[�e�-;*�����_x�����j&Z����rs��r��������=4�+�=w���?D0n�+���N��/{H��e�P�&p�s"��^���6�w���@;p]�Yz%�\�u���mNJJ��H�N�B�����g�E"Q�X7_L�,dV��3lhA��ѻ �zE{>i�m�����e��f��Έ��B���G3�焥s��r�"��@C�8��l�G��ߡ���������U��)�>�vO�:���)Z��?�YB�p@;31Aȩd�TU�`����Y�G�2�!�_�?\d�c���:ʝ�,��۠��g�e�M�R�xp�@�V�� =���*HD(a,�FL�i5�g��i�}��K��W��dSA����08�~��ﯲ����Zt���@h��6�N3R�մsҗph�����./Y������0ZkU��9�3a�w��n6�V��r�GY_��¶ir͋5�:C���KA,�6§��L{�r�.�Kk�~MЅ�`:h�H9E���T��Í'ؖLK96S� ���L�B_	�"$^���=�o����ɣ,ZMY
>j�n���c�ncȍ��]k2���Kp�{82f�wa���;����Ų���s��_��ie10�0�7IN�]!�6W΁5�
�
�~��͕��Q�´��t�N��e�X}?�=8c?�*||Q~O��j z��k��d��!C�+<ڿ����QB;F��-�wJ�68T�a
�_nvvsb��7W:���Hߐp��=��_;=��~�H�:��=���,[���2$wbY����շiap�@^�0�����Ɖ��X�6u�����y��<��I�Ex�v���.P��ѣ����Շ+L���'5����>�\L��_���k�� ��D��`��t�Du#F�G�NV�P���()�LW��d��M��rPa��mL�H�9�Fd�esٖ��\�KѬ.��׋C���L