XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���
R\��&`#3�9l�߾=��C=#����cE�v�!:y1�)�źH�ڇ;���6N��4����2sף&պxU9�	�eX{���$ݪ��=��ғ]e��8^�\���C�6�������)z��b��$u�
H)ЪI�i4���o�C�
�T.L]=����lZ��&O28��O
����$l���ֈ���}�$��Ʃ鼼^������O6���鷞�k�h{FT�-����n��@NXC�Ю>^U�Ra15��%��B�wttl�2�.��r���e8֔�X��Cb����Q�9�<���6Hrc�6��K��\�6�]®�IfEn���*� SWƅ*� �:'CJ�'L��Mjcڈ�W�Y��u�YꔍQ+|�����}��D-K�ܟ�����J _1���Q�4S^�����7<T���G���M6�n��Ba�_�G;��!�<#\C�֢{!�t����oj�;Y�oϼ��S�} �p�z���y�5W�s��=	�-��R��<qH�5�~���J��9�ٶ�KJ�W#����qLЭ�H���V��ԕ��{� �
��L�û�aS���^�/WEsd���c��y���I������RMN�>OEvK0��;N`��7�pV�P��h�rG�|%���xN�K;��K��T�O�����;	�F���h���o͂:�j�|����6���]�I4<������q����'�X<���Rj�q_fSx5�+Pݻ�/�\2UQ�d����u��_���(���D#�]XlxVHYEB    7744    1780��uk�w`D�J=��ez+L�+1�i(_���j"(Lg�f36.X1� �O�}W����+����#W�h�گ^� ��Hd�����IW�_�W7�./{F�Ǡv��#T1['2�W�R�[�0�6���p/�y��{��$�`7���8�O��2�Z��F��<'�5��D�
�m}Y�����:��e���h�Ԧ.��+��=�q �h+k��WhK���hrP�:@ۤ�%f��Jb�	�H��Q�2}G;ϊ0����NcR�!��ۼ6ho�m[!IeaF؏?j��%����V�sH�:��E�woqZ�9���[�7rkrtG�.c�����#		*I����?d;�f+×���������(a; ��L�Ib�`�nh��y�mf�&	���P��u�ϗ��y�㷐2��58=�8�E�(nup�"EѯRE��<wd@G	@BF��?��V�%�c5��If�d�!ݼ�pef�����#��,
�?��4^�wPSAK��s}�����i�r�`2	��C�F����Ѝr훊���@eџZ>�^�
@�;5�|YZz�ɰ�k�0�g�,�L�VD�?��͎Wv3r~`k���G~7�����O�6�ܧ,��w�'���dW&d��`�"\��Y
�<�ٝ��b�B���eH�f[t����m��l�P�eE���G�?�=!�v3F����
5����w��x����XeÍ�}+�6߹��U�VE�Mi��	�t��^�}���6�~��6kQ$[�pBW*��W�6��Q>6��F����
=�j��(����LPKmdN�B�>���o,���2������0�3y�ON�i��>Y�+�i��a<Ɯ$
^�
����R��(�������jv�W��;�.�
\�<�jD,z瀯�$��_1���&U˵7+���L��5�3��D�6��e5o�2_.�*�D_N�e���K-^\���e(9C�<"�E�j*�ax0fkl�
޾��O$P�)4�[G,"��g�RES}ZoUhק�ߙ 6&��i�%��� �,��i?�\+LǑ}9�p�\������yj�q�p�tU�<��� �zç�����[������[��ڮ��y�V�l�"Peo$���*��ku�
s�'	�ҚX�1ի�
���@m�UaߥQ�ةʪֳ�ώ-1'��f�m�_a�� �N��@��z������W�V�* �l�=h҇�)������l�ל��b����El�_��݀�D� ��KV�5>�P��������R�n��~��c���0
j�X0M��*����M[�t��)���)�:���ĕ�y㈆����Re�,>��7��3 �^L���0���GIF��{�<�@��%�$8��֏!��Gu��2h��L�K025��4�͍�x�{ x��#�9����������y���7D�_��4!��h���5�M��	�ՉD�'�)�P�|ߡd;�R@�V8�&Q<l��'#�w�E�>}���v�Q�G�q�=,�K�Nc��L��K�k��<�N�Ub��on��E�!���&'����$��K��[�0�=��u�fk�b)�j�Ynv{��ѬXqex\y}|$�OO���@(5c��m;��La�2M�n�������(>8W �+�@_��n�2?�ٌ�бm���G]�\�l����(Y�|���0&��Ƽ'R�4���j8~c�hn�7�~ �u��9��[�Cp�|�� 8����K�@4ʹ_mi�x儆D��7���<�L��A��2D�䨵�[���,y�E��/z�a5����r�l���R�>@��7��x���̂�_�OlRjHh+L����RYF>�Ɵ!s��V�2�f��}
�$,wa�F�m����]%a�������w"�Ba��&�cm��#�F� x�����av������.� �?�Y���`�H_B�dZ��v�hA,�5��7qj��g�R�����Z�Z���ֵ���0	r�a���xyto=<k���#BGr}!	�-O����%��Wf�VVaIc��A�-$1+*����=J�_yΘ<�ި�=_�5y�~v�����P�u���<��N*�1R�r�����3a���DxOi���I�M將�1��17Y]:����ۡ.y�4|c_H<$:�D;6+`�S���v�V���P�\·)B{��	����¥���Д5K�
���L\��G� w�fi�DW Q
��鈰�1��3�5�X�!�i��L�]�/�N6��ψ	AF�1V!Hj>ː0� &��%/a����Ѷ���� ��ͳ����k�+T(�7�z�ˆ�X��Lk�� ҽ��,�(���S"�D{OZ]���G;��!���:
ۑ�Qh�79���E�p�Q#�|e��!����b/m,����R���E@�G��|�2�i2։}^�9�`��Y����"t6�V�ף�wh�nRMy?�P�Y�a�2wuP��*ػ�\�xdN�ӤU��b#w�=�]�|�|�D�>�Y{�~b8��a�U���?�p}Lh�l�|�����&�Uٗ�|{��Qis	f.+k�A0�!��0G1�{��Q���p���+�	�L�5�T�=�=9
N�T��(�#9��;T�%�q��u��A��*/�N�\��j�!\O�vqڷ�f��d�g����z�����N9�ܯ{�b  j�Zl�O�(�P<I���-��P/Z���2(J�͐<�u�r�?����
!S��*��N#�G��n�������V2ކ}���UnI�xTZ�C��c�!H�j�Ό+w�?̭1�%&
���q�:���V�J\�*zT2�-��X\��Q�F�*���Yh��C-+���1�l�1>�{u��ґ��(�����n��l���#,�Hf5����L��-/���ØD5��2�9K��<�]��@��b�^FRG��ZG��s��2vjv�df�e&�q�ɒ��ߜ㳳J��P$W�^h��a
���?�].�~T�1�� �=i3�-˷6R�|b�N�U��ir���5Tsf��W���^�۰��&k�э�W���{=@;=�$�>�W�xa��O5��L>�.��m�izt�uȒ�Q�+D�X,HD�{��?�"�7k[������ �,�oj�j���+�}`r�����qZ4r6��F��M�_�+�M�H9���P=E�mJ g��*&����O��J��e@��R2Y���-A�I���b ��<_;�)��Qs�KǪ�o����mV���,��v7?���d�,i,���wm���kD��/��8�
1^z�>T&�}!�G*]�	�vc]�~��IGx���h�-�s�\�RY��/U��A��v�����b�ԩ'p��Ѳ�8����x�'�Ә�B�FMPQL55�JB�>�5�X��K�3�3#a"�Yt� 5dc��RgJ5뗩�	���!�Em�U��j�>Sד��I��鯬��@o�Jè�>���q#�]��d��̹��¨��ګ�]Ѧ�m���Oy���٥�[�U��6��Mj=
�:�_x=�:M,7'2��&�z���U�\!I�ׇNC�~��{��6qb�a�Ŵ��,�ڄ�k*���]�������Nc-��� �0a�+���'��3�5g�)���";Խ�ꛅ( ����oQ�f����TB)�q+�E��)Id4#Y̚�n�4X��pUbV�T})��S�"Ǝ�}�%����* �?�Ͼ������8�G�C���<��Y�}��W���޳�|����Da�*Է�g�y��������?�+�9�߬�����L��&����.#�b�ys\4�\�n�l9����׌�7��G	��5���/�d�+�C1Z��qD8M~hw"ňr�9�_�9uְ��������*ՔX�yU� �>���;ɦ�=�����H�{�A3�̂V��q0!�ͱm�X11���{1G��z���������H�et͡��;VN�]�H��T�4d��0B~e{�M�F�>�w�����*����vf�Ϝ+�U��QϗK��v���C*8Dv�/�5M�K��d�;�Spp0��8�&��w�m!n"���BE�B[�C$|!!�6�(������:|g\c�@�������Q�o:Q.�j��A+j}XϘ1��%E��ɤg���#�)��)���(�|�n��q�NxL��#�!���Sj�t ��||�(H�2�>n>�f���a/������՛E�r�8���	H��y,�N��*�@�bh�.�"�f��sѓ}����{㮟����hoYefdhgm¢$G�\^�͊ah�y5���;_XW�9�z<���m�����`q����n׼v�&�������u���p��6��A�Q���+W�7��p��t���+�� �乲ݕQ�9��I�N�R�����`��{�)��,��M���q,�<�ց�~吡��u�h��[��R�pr�nV��R������a���j�crcIT�� ){��B��\�?���&� �	l|��b��T��T1��U�4W�E��w���f��e�F�T��xaI#��L^�L �,��r53�hT)�h�R�5Ҩ�$�s`�F���D�dS�%�և�S4pq��*����z�k�i�G��j�f�/�K��	� �'���~���{�c�Ie�!��>�s��ؑ�|}k�6!͒-Z�?���1Q��V-IuiE��L�/ ��}*&��>���{�����M���H<�x�o	<��H#%�by���E�K\� �|/['hk�ȼ�/[)D�l�-�
\��8km��S`!�@>E�PD=$}�����Y�q�ե�v/���BO���Щ��<��X�h�i%����_�c�x�\�o���=�`����8 \��aW�>Xl%v;���[ڎ���/��#�I�5�r�7,k�MhRW#Ď�Zֆ�k� ���h�&��:�pE?Gu[@���}�!P�6�������!�f�3_�6��@��ᳯ*������n���f[�l�B��9��*��B���?�'�i�u���ڠTi���k*�G7ڄ$Ur��Z-��/��>�W�ƪ|��vU�<�|?��d'�j������}�Jau�=��$,��<!����f�5��J�J�d5@�4G�t����kC�ɶ��A����!C�i��k���O5:��t�T�Y�����ӳw}*�0m~���|1*.���$Gs�ш:�#�n.h0���س,�������Rz5)��rx�GzP�e�ePW�4s�.���q<�[�ܱ&�Vhc!�1Rr29QT�'�Pp�S�ʌ╶�O͕Ԋ�E#Nĸ����;v�cGH��ȵ��w�ZV\9�� �%긥DZ�4�_s󳠸���$0M.P")<�� �2��Zՙg�q�p��r���B����I_�e�ݔ�|�E��lؕt���fC��07�h_Z�S��pۡ�)^�1Em�N�p�$@�n���.d^/��_�����^��)w�������4�xd˞Rgŷ���X�<��ڻ�U������ٞ&ߣ�!{�)�>PJ1�X)0��+�9�h����!��:W5�1>�<=�q��p�I��1힜=��O�-�NO�iãƱJ7�=�ų�M������3k������ǆ�T�]N���t�̸�"|p�x�
����+����!z��:�	t��N���p�I�A����?@���sx�aR��Y����^�5�H�m̓c�W�[zt4˻w�f��a[0�A��
m��S�569H�������u��8
�D)���K�H㊾UQ7��m�����_�`����3`$X`�E���l��{BB���]饸�;_���nY�a�n�rؑ�g
��|v�?�&���keq�*L!��nK�����Y@����ĈU���e��