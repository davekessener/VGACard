XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L�X���˸
S؞4;������s�y�o�=RT��� '4�e�Ds�ʐ0���ޞ�9�k�{&k��dv�㿟`H��	�Fbv�{�n.�!� �h�XF#�zu&NP�/ͭtdO�Q����Zt4Q�1�{�ғRbRe#��0XHD_�F*���X�����B
�-?ت�'R݆6�̅<x��L#=w�>\��suۼ�$o��o1,�?��y!N��Yx�������DN�_S�q�E��@Mf�����[E�����z�r� 19�D/�����&<N��{�����%�z�����c�p���lD\�r+�.�M�}�Յq�x��F�������1
��{$N�'�*uZ��V[���H��T�6L+�jکf"e���L`��G�̲��6�����c�WJRP�]Z7���.��d緁���$��VjC-u<_i8�K"��.�s�~0+�{¶z�}N�Mu3h(�Z� i̬�	�f9��S#oh��tj=-9(��K��3�/�>�j�����F��[�SZ븒).�-j���f&��D��_�m$l�N��At�eL���b&������4:mpb���4U�{�Q�(�s�%��.�ق�T`&�PyZ��Җ��H���x4�������M�B�r^��K	ool��U����"�	�.o8�Y���K���ӆ��д!�3�?PU��2�9�-�hW�'Ể���_�l�2=o�dUDR��2[�*��Fj�Af��?G��?�?|�E���ޣ8����C�XlxVHYEB    fa00    25609�r�5B�]%"W��fdi"���$���e�qL�����W��]H�w���
��R���A�@]�K�s�A�5(&ק���>�KI�p@^��MDP���H	 ��T�~���3���!6 �I����a���u&�H�0���tӢ�B�7�Y19�&�Ũٺ�u�����+������� E�?=C�Ȳ�5dV�dð��T'�	��tv6��t�ԑ_���6yxѕ��@9VV(���ߔ��a��j��nVS��(G�D��I�]1j�.��a6i6R�vC��U��2�
��쏅��R`�U���W+s�́ñ��Z�ͧ8���P.�A��I���K	-r�Qb����t�1­���8 ����pip��!���4(�!�f��a�(��r��n�8��-m8< �΁�VǏ��<���c�����ښ繕�dT�����B�:Ք1}�j��'P���'��'�G����_�G�C�R�p�I�#@��)%ɩ���2_�b;2���O�]�춘*��u{)���轩3E΂$Dt]�;���+��4��M���i�1aci�Hr��&Q�~��C��WM<��J\�� ������Kj�-��V�������lۙcS�+��l�aoq���G:�`{
�P�hx�Ψ����Rt5��GeH �$��;I8�j�D��;�[aT&*��,�<iV��7�a�H�m쉦�Z	t�����Q�l����-E�G��Qw�A���@DϜ�ƍ��w�_��-�;r��g0� ��I��"��x���,1.�+b�P��ٖ��^XE�C�֔�+�����hL0�#΍>Rhhi�5c+�*�+9Oӳ(��gf1�^v����Ǌl�Т\�z�S�V��
j��31?��?��z3a�j����ò*0� m�����q��bxc��(��HV�����ٴ�zͷ�06S��9�5 a�*�U��-��Ss'V�s���z�
I��M�E9�Kt�-��/���gw_,�]n� ��7V1��m�"=!!����Q6�`��c3�6��R=�JL�3�ʓGEͪ]��O��\6��mk��:�A�d	�)1A��ߢ�1�еWƵ-�`�Xdz=��|��dN�����<��K���fs�,��J��k��?�a���lW����;iYt`�社�o2mcs2RA��xi"��3��e�9{�o9�[�� �	7�Q���q�؏Ċl��0fdk�c��44�9�\�}�a�&M��_
�l#R�Z��bv�o�rQe��uo �S7~�~�N0��W�����+�#����қ��e������Rg�<�pR�1�V�T���C���Yr6��@p%�"CZ>�U����#���͌x!U��=f"w������pf��,o�bW���H:��3(u&����� 5��a��"�3���_Wl�gXy1p��%�Y����X~-~���C�����8="�k���֖��(.?z+��,�˴��Κ��[�sP��H%M(����j��^`<�{�Ɖ˅2�����{�E�(s���X�(J&ĞZ�����q�����W;���D(�@R�<p�T���M�@O<L�����Um�Q���r����~ ޹�3�Ve�-�0�T�>�������ow��6b	Ӆ�t�'���$�7�		��*j+ĝ���z�¤��2 ?6〡�K��=1yMvƬf�A4ߔ �\>q2��U�e)�Ż��ԙ�/��lA�q�m����7D��\3��y�j^��>���(�(�f'<�fݱ���E��7��Y+�caî�߂�BN���'DF��T0����q�D���&_E�~� >`��x�st��$6��0��:e]|DwZ��<�w�h���~��߮!) ����
f�R��d.mT]�A�	v�i���eם�孎����xweI,X��h�[�r�ʑ{3"u��K�F~!�9�rO��~+)��
G�M���|6��+wGcϒA�7Q�}���G�M�g9�A�	�Zʎ�{��+�>����E^<}��rg�ۻr��48��=���]�O�!���-�ڂrYv뷹�s�B"m��"]�q�s^y_���5�Җ��05�^C�5ۼ��	�:㛱���t�e!��VL0��C\�F&���Z�w����<��mu> G3��I�+�M���$@�]�?[c[@L��I�y`upv�`�����R��w�~��TPP/��b0�o̩,T~��d�T���G�R��a.���%�H3�^���E [c���8�J�ӄ��K�/��O�|��	}� 3!�d�+�s=g!D�>�R1���z��@]�Ty]+a���(��Myu9#N���Hv�����3�9
6�������7��y	)�C�6���-�n���犘B�!��R��ho����W���� ��ʦ���,rQŏ�{4�5b\ﵖ`
�Q"9sO?���엋���t&s��J��������Ί��mv�&#�6�%���m�H�!7w}�-���H�^wI����ٿe��F'��6`��o�&�t�iu_̩c�~��<�`�(�a����C�a8�T�ѷ �s����Flv)5u���t�C>T�\��!�\��˾��&�3\'ؒg+cQ�7�Q������LP���b��ȊW��P�O��m'#����>��z���͙/����}1�}'M8e1����dx��Y��p�����[W�� V��D�u��}�b�0xC
�)�wb�?� +��і
��R�����O��|$�K�E"d��S)C���[B�vh
�ې�H�%ƅF�ݟ��_�K��bؐwmbn�}�1��m��X�I�]��N ���1:���������-�~�^,�����	e����"�x����ᒣ�Mw���L������?�����:��)�h�j(�-dyT*��{�}���d +g�ƮT`�g�_;�B�eA�77�V�M�l�b^�C�2���ϲ�k`���IjY9Y���
1�\�����'"=E�`G	o�n�_�Y�g��Al-��45=ÿ;������x`F&\+ $��gq��&��05�	��mw3��?����!f� М��B��=T��e�#��]?���e�H�I0=U��\hv���h���+�K��i��)<a~<#L���>�/\���W$sQ:4�ܼ���h]r�)L/��hI��s�o,��'�#7$���O(����;ι&�L���̰��n$�ت?!t�禇�Q~C�˟���NČyv����W�9
��V����`��f�}�q}�?>��N.��h��������SK�Jv�sE�V�8�TS=AJx�31kw�a��r%�*��U��vL�$ ���l�>>(�H*��ZzR+Է�n�;�s� ҥ�38K�8����Ø_z#��El�������f���8�e/�9��!g���(G%7?�9q��px���;m}�Zv�Р&�.-��h[����H[tB��Roc���.��Z�z�����_,�nx�i�O�뿁�Iksp�I]��1YS��##�~�Px�%���=}�^��9C�C��v�H�#4c�^�mwD���x��R���]�;�־���6s��s��V��աa���_���q`,M�� �ך=�V��2�I�6jxƛ����5I��(]��t�{�ഢSg��;g�I`2e�\"��� �
����g&T���g�t����0Ĝ@�_l�{ufl�}P���!���K&�p	���/��30)�d� +���ɕ��[im�R#3�aOڜ�4���ԕ�v%O���}lw��1�U2�g尬�T9h�R.)7\�*�8��&OR����2�]k�;����J�z��rZ�� ���햬��ܔ�7�1L�I∂������~���)�!�Ҿ���( �ߕe�[���)S��pP��Cs�v`u���3�ꝁW��_�g�fv�0���=��C ��>�K&��V�6���ˀWXB�C[��$�x�6�ː]�"v��4��ڝC ���[��i�5ΐ�C�S�*@�	�o�2�`� М�ۖ��Q�I���~���}¾ �� NR4.�/��}��h7��K��
�H5���e����'�G3|��*���e)t��nF��!�� "�u�?T���׽{_���@���!Y,B?ȶ��盂8��Kv%k�@A��V&��"�ɗEn+�P&�
q2� ה��8����c��8cn�jE���ym���� ����6+�)�,ܾ6��K�&3Հ`��$,�}��F��:��6o�f���sV��Uu1 `���a}S�d�eZ93{��K�~�w�R�L����|%>�A1��g+�s�	�r���w��۠���O1���,3͍�>Nց!J<�,e��Hk���g�rZc���@����R���6���9Pa�Q��������s~D�x�N5��bK�I��˦��.�WK,!֒�8��o������Iཡ����xG���XH9�W���F�U�����S��ŋ�J(sN���ɻ ��"a'��rݒ�  Kr�Ľ��&C���a�M�R�6s�b'~Ml{b��c��p�����8ɫ���ѧ�g���-]}��.�ʴ�����=�й���7�֕�Ww�]]���������y��F�J��L�Ѩ��$u�/7��*Э��C��� ��4S�J�'8�L�b�x�Ҕ�v`3��<o�Xe.�� c- q�ޓEd��\�~M���u|�	�g���D���4.q`�1�߉]���0�xzC�pGBx����^�/��5_���PX��)�������Ƽ�/� ��x~Ay���T��敖��z=��x}s��]�ߞ�{"��lG������>�.lJfz�^(��l;>F�J
�Ƌ`�&�� �(wW�	�u�a��?�pH����P�Oj��!����-��k\��1f�k��z�� ?�=�}EP��P�.�&�97��J��3. �43��Z���ط:���#�'b�C�]6���[rT�cc�"�?�i�I���iș����&���f�w#g/+6����T����_���_����_�;ib7�P�=��^��� 1�_�������ْb��}�6MU
�n�}=Y�Fs�ѓ����뇣eh�cwCt��D�s���Y��� n.���]�w�����%��`Í`��p�]y�N�l1{��<)� =���<�ĻL7��㣶���������vk��|�6�UP|6̂�s�U+��+�PG#Rsj`a�6z(��R���F��ei܀ 4�dq����Q��K6�A#�%����?`7:���rt�p=�R����>�tt��8�F�}��W��	�`����l�	�k��u6����?�x4\�ʥtFL�W#�~���l|J�ᵄKJ�퉴��!��@��q����=��#����_K*��E�TٝE�#�����d��8�_~�)m���9��JA�ų�I�<|��A��'B�?&���rk���RRR��L�D����9�Pr�饺=���k஬�v��o�I�V���
���jV�?����̐ ���jz�J�D������oJ��g��Q�}?�mҔ}��;qNG��\��WD&�,�4��xP��t�I���q9.ձ����hGt��zLn��>w��R�ɓ�Yt㞷~]���}Q,ؕn�K9o��̂f�%����ct"�8��<���`���EM�s���3��9;�G{4�\^�hJ�mp��-d��=�����d�7�7"2l &�����ŭpMZjۜ]���:��Z��"!� ���_p���Ln:s�@\u������+�C�u���֝O�LY���tF���[}�����C�]��IR�$�D:E�#^�f8��(��>���1u�xE�	���jk��n�gw�\�Ob*ґ�^��Ʉ�)�����D����)c�-���������c�O�WA�C FU�
��<"C^�*�|G�7Ebr�Pt�Ҝfo���&Ed�C��� �_(G���ޔ^yn��K�V���aL��փ�|��v� 
3�T�������o9+���U7KN&r���^&�1�avtɴ��|F�O��lz�pM`Un��D ��+e����� !̜��}�Z��������w�uW�߲I��e�-�Ϝu����,ա4w!H�J��a}<J	 ����v��� �C'�
J�#��P��NR�HwŪ�m��;�9���;���A-w��pOKTB�V�J�� ���?�z���v6�����&ypt3&9<�L�b��+����C>��Zs
B")>Oo��e�����"Afi�04��c	�(�ڡzi���� Q?`~\��~�,*����Q��eEn��-h���8��I�	�l��Vs��{�����n�����7�CN?4�}u�W"�E>��Z
�Ν�������!L}���"�J�o�I�6H�]�l^�� "KJBC�l���OL\4��K�	�Dn��=T6�jRG��=s�.���X��[�ňoG`�[�r��ZY��a$S��[v�=r�Y�l�����Ր��Z}FZ�����+6\�<��ı1%��G�� ��5��r�qQ�����Q��G;�K2nҲ\H���>ۢ�0���	T�r�p���=K�������):֔���M�(�:м0� ;<�2 S� A�1|��S]��E�cZ.7^�U)%�4*NCs�hR�؀4G�|���a��N��!�K�#Tc)�"�jz����laɠ�Y\�I��}Y,��k},F��V�}�n��1�{��xO���SA��(�~��}����,�d4u"j�Kr*�6�J2�R��0���f@�ٸ�`������v<؎p}���qݸqrV�!��I�p�BZ:�����wC>�ѷ�͚��@��͊�L�/ Ҝ!]���u߹4۬������<6�ND�@������0�'����O$'��c��1Kk}�8��j���aF�X�N",JA����������8R��8��ޞٻ��$�`IH�#%�d��&4=Ŋ�B~A��R�~{gJ�|�3���p ��Ti��%/$
<�ѣ�XUR��Ɗif��7ur?w��y��x��w� �6ہ{-6�ƨ��8�;��G�C�O����]'�X4�
�brF���r�'�-?���]��]��}t��D����	h����ٜn#�.6�/�!���{6�{1�3���{��79���7Lm�B�=Bv�������e,��2=�7/��x�8���Y.����lz����K�����]<
��r��HO�E9R���L~{�ɱk�m����Q��'J�ݾ�2/��}����}Q���V�����xzx�b�R��|�~���
{�P�,����N������ؙ�FX�.�<�˹��K��H�đ��L��K�f���#Y�ˡEG�P(;^ͣb%*F�������A[K�q�u�zo"2�f,�����Ryc�O�;%�k(�R��{"wS�|��S�B�>��@��>���ќ�7���b�Mv2��p��J�I��o�Çڥ>��i�{^������>j���W�N����2k����)��0��P�Y���<� �x�٫�	�}��}c�����R��f�M��li̇89��������/d�˕3Ó�x���H6E���E��_W�b������u��sP}�p,AR��x�`̇�R��2̑M.C!�g�G��̽A{U\C����[����\�&���߅5Օ)/��T�{��X���(Kc��s Y���J��s��Q�/e:蓑���`��ѵX�����ny�}�/9�װl���[����a.\z����~�Guz���R���}�n�b�d�X:?8��(O�l�u�����m��ܻm�YU�7��ըFke�EK3�^�-k�uKz�.U6����U�/�����] ޹l���7�z��
����BOId�y-3���n�7÷={+h��+��!��[�Y�����B��NU���[��Jk����k���q&f]�Jf�NOM�[.1��}�C!5�U���+��d�D��?�5u��:��A��sQ�����`����"5�`�3�EJ���,`��O:� J��J��Q\t!DOO��_q~�r�s��<*�j����W��Ê������4�	/$2��# ����U�J��NW7��+�. Yշ�9R*|��Ti�/�+	L%��K����l�0�m6�w }'�ɢLL�����hx۫w�����$�!���KX�-��F��]4a�����žy=�PL��;X��%�z(��>8К����*�nfg)�/fn�c�!��<���lTvZ:s�g�>2��w�9�������'�;̑):m�27\0��9i�4��B�@l��ަ.�M6b?���/��e��	ͩ	Ư��y&L�����8�	f(/�_06�y������# ��~NӶMVG_YQ��8e6?x|�3#H��I��ެp���r3#y=��(�n�Ja��AlWK�UKzA�Oܔ�V�΅i���*&ݭ2�XӅ��-q��K��C)�4p�5UwŌ�L�n�BXĽ�[%�<H�D�R��Y�Ew���^�m�y[����!���$��H�f׸��g�V�*\���'��]� ��ռ��V}7ζz8?{z����B����0����/u��&]D�#���d&dY��``���Bm�{bp�%s�71^6{Y�7�b~	�&���2����f�?��jm�a.�9�`��FS�sQ�=ڵd�U�+��jʇ��]��#lV5X�e?��	�� ������G��fC�/��m|�$z�*�=����@�jW�������f��{���!���x!R]\�/��P��y��?Ҧ��E�/ �8G�ƃ��j��z�?`�����1n;�9�A��@?��줫���B*|�d��}�P�]�_)���&2w�����o��f`�Z�,_��EH�(��tY����&��z�X�>���e�j��G\�S����1e����d�T�n�ދg|B�EC)�"�B����=R�/�"��_>�Y�ht�CWy�2�	�)�H"�/%��iQVU�� X��Y�\h�N9�-(�L�=d�.i�n�J`XWf�4�Y����c��_X��,����Y���	+�$���yk-i����`�����8'����HZ}�Q���xY��o�xx��kH��_��֝��Bk�H��*��@���H��iz(����p]�++s�o=FE�+vO <�:���a++��怡�dPN�@g���+5��	��4@���X�����.��+�aSA��Z"�OU��u��Jv�%A�c�*�����-P�{�ƅ����d���1M�\r�8�H��"]�h��$�X�Ƒ�YXlxVHYEB    fa00    14b0b#Gݧ�>��� RС�U6vL�jB�hýOL�s7��(����-K�I��g@�2���`V���:;[>w�	!��'o���W5���'+k r�0D7-������u�`�ȋ_q��Bڭ�]�
�$S|�5Z4S��"=�f#)��t�Y�����h�voL@���V%���P�%�qf~B,�����ꃘF|��c��p$�4K&����.�j�bf�����ˈ9qu���d���>d�ӾV,q��w���z�������ẎQ���[Z�F�J�[RA�x�k��P�y.�9�نs���w%��_�n�`�����j�OO�q�9�@J����WP��R��e�)�Rd�2�Ja�J��l`ȴ�3
��\�EA���N���#8��-�
P�Dۓ�U�/�}w���`������/������dF	$��f�YkC���׾n�4�Wsbc0�%cٍ�@�P.�r@�1lD�.6q(��4Q���\�@I���&���&U#��#|O5z�Wu�t�[��tc�����a�H����"L�b���T��_��� ��CA�hT\��>�rQ2N�56w��~�6�yB�1�l�.��:W�v�U7���!��h�9pb��(��O�e!V�F��󃠷����:>��p�U<��tǡ.D��l0�J7��+�y��˰�K��OՉ��1�-��&���0Amf�����(#�'I�M=�Ĝ�����͡����_Cǂ3�����)W3�O�:���	�'ٴ�?PPw��!-�AS-�>��1 �:P ��Z�|����R*�V���k@�z0v�p�K��b����N��p��n���[��ҫ�t�`C���M0��2�aA�[�� ��ȆI�u`׹�����XF���]!l�&m�U�2�f�ǂ��K���G1�=�b�et*�N�m`�����ld�?}���E�9�^9��%b�°���:�I6�iZ������=��D���+�3!�� �5#&��cL@������ޓ-6VL˾�]jǶ<����J���ޛ�0��g�����!�ԃ*df��Ȣvs���9ʎ!݀֖�ٹ� ��Jz�?4=c�k���rM��Ѥ[�q ��N���Q�� K�e�$	���s��6B�:uh��j�l|��eꝪ��y�]%0��)�Tb��g���Cԍ��U3=���Y��x�>*��9_g�t~Y,���QrL��ѫ�iנ���06����~�H3gނG�i�<LV�R�8%ڤ��GZ���`o�X���V�:���`��B{�#S3�������׍���R�ݳi�g%��.v�n�_�Bq�.$j�k@�o�5P��8ѧ�S9B�D��Ÿ������e�Kb.��]�8�}4�1�s�ۉ�A�����g�R�X^Ko�0X�Ľ;�"��#�;���mLy�;�J�ͻۍ��$����U�R/�}R1!�����I%�-�f)́!��W�O��u̎�uHl�n���x�cN.�M5�b�X��jȺ��Ulz?��Q��t�1�]t]-�"ᇤ��>�"�߉���	���p���X�wh���9�H+km`wK?���� ���T=~5���\$'��H�c���C�ٜ�+�7�4¯��In|�j�U�h?�������O������v|6}�1&�cw�0�:�ZE: Yz�+�{s�S��f#rBζ�q*�*Wv�zߥ���g"ŭ]\%�^�6����IR�f�rߞ �q(q�T��*��ƺ˞�?�4��#H���F��Ch�aj
�ZT'6?0�b�o(}���tۂ�:>��ddIa�6ƥ'�}>Pa����$�v���[&�	��1�$��	k����2��Hl�d�����i<l�,��ӳQ���F� �cm�,�>�~��?d/	<��鞐��*��\
}�T�0�T���-
Ymt�!�6�z��}�QK��VV�*	Mߒ0�q ��Q�.^��O�����;!�{YP���?���Y)ݭ��ȷ�wg��V�3���C�rY�T�/������h�[R����,^\��~(Е��3w�?r�'�}�=�������&�����T���w�E�V�H- ��9��ȪүŠ���K�m��8�q���8u��})YgU�=�5b�:/L��D��Z�jO����c��E@qP�~`�����o�g���cq7es���t�Ud�5�~޹���<�iWj>+�璖D�̻����������ћ���a�s���ͦ���w�	}�)��^��7]�A��Elw����Tx���˝�b1'�p���ƺ޼�┗����f8c\d�Д���|���!&�����ǋ�x�x�[tj�"�h��e@S}2�C���)<*�Y=XJ�J[ ��5�Ö�֚�P�$ٟ8I�_H2i �����i[s�9!��-�	��+���!9^�4f��F"��-8t�\l�A䃹�4;��+ձ��$����O�����[:0�R�]��v�n�BI��:+>�o�g��z�o��u�5)��>��֯���}�|�2e�3�K�ٰ��R۾e��?9�&`�(�-.�6�@(�\	���V$��S��27X �Wm�:��S���j/��cr�6f�J�gG1uP�S����?�t84*n��D~01�27A�)�wR�Ǩ%|��dSVt*��3�8y���E#�F(ǐ���6�uA�HI��Y'���Z�ӫ�#�t��\��	9�1�Q�%��T:*�OY8�c<T5H[�����- +��VK���=?@J���ƬoYϪ���iX]{�;<	� XcL���
d�%��tf�QG�\j��|Y�꩔E�ŝ�Lx��ȅഐ�h�ͪN��s!nCu=�C, i���լ,���)h�*F>k���`����G�(��	�%�d"oi�CpZ��g��"��\��`W@a�0�{�����x�W�+Z�b�ޱ0QIs�u�{q�Kwp��T�˾�;�T���*O��al-#����c�ٜ}���A9��N\���|ɑ������p��g|����ǻg�����.�\�!�4���7��nT���]�/��&�����I6��K��ZU�6w�ȿ�Rn���o$�x!��_�~�7�u|B.���eg-��������b݌оl��$������`����RF�H�p"�s�o�
w�y �� ���fp�Th�s��(�-s��	
Ԥ�Z�R�嬻��w}F��*��T�|9���ƛ������⩸���ӽQv�������YA�+_�Er�3r�Y�l�w�%�������)�,��IC�a�\��~��lIq�|I�:+��O�:(�n�����&Z�{�o,j$;dK�A�f<.IDv�֏|�.*Qi7%��7k�Y�Ĥɽ���UtoM���aۃ1���scl��
�R��w�Ed�����g��`�	%]E�9��#qu�&�ʤ�R�;c��;�WS,:(F����C���%���Ɨ*����j]4D�´#��j��5�B����7�/�^p[>����M@����+Gd��y�ܭ-�67Qem������ˆ�#���4�/K�?������*��8o��'�=9���<�	J�,�n�
R#���@�h���ʓ&�
��o6S�Pw*� ���i��0P�+�����F�)Kd�� ��v��Q����D;�]/�]nR�$�!4��1�R� �c	��șS�x�m"�8,[&WDI���)��d���[7�bj�n��Fa���?�X��9��jj|#=��n����o�]�E��I�F�U�S��p�ov��0ꛣ[�SN��P�?*�ȢJ�X1\?�+���x��� �b���X�̨9��C#���p/�걄ȟ.�w�+��[}����_���a���[4N3�7�ۘ�_��8�	�B^�n���S��3c[����n�ǟz\a�9��XlA=��u��#�؁�y!�R�-Td�s˘*h�Y�RM���|�Z�_uR� � |�by�]�p���Ƚ*ʪ��G�Ы�X��0��]�����h����7��22���[��%s�a�����k-?p��Z��
G�ȍV�wB�Qd���n� ��Hr��������z��*��$F�	"�a圩c��(Ѫ�	�m˖�=����~��0�B����ޅ�s)��^�Y�t�����Yf���̍rO,�5Kˎ4WR��f���u&!��@�߫Vn�X!'�!�E�tZl2&3[���=�[S�|qOd���@(,c�������Bv��Z҇6N�^�a	�0��5ڶ�E-��k<"��� ��v�~/��U�Ҹ��Gf�B,X)��Κ�=�C�Yٕ�g�H��
��7�ռ��Q�%��Ֆ�(w��l=�z�'���=X�T#pM/Ūz�1`L\I����_Е���E�γ�d��ʹ���33*|�):;�zY�i�0��!v�������&�"�����4��{7	��E�\�%��y}��W����p���T]'�K�4}b�p�h1���+�4l䢙����t��;� �,/����0e��KM�p����=��x�3i��a�5=��nβ6��>��5s}����^�I���vS�6�eԆ�ʒۚo�;o;G�Q����� V�I��|��N��B�X�C%w�۱e?2l;�	ɤZ�Aі��a`����2���?�bE��f^���@tz�V�k�����?|6xp��J��ym"h�YΦ�y�TX!sj��z�x}�r<�\�t�t,��x�D啛����PQ��IS���
���uZ�V�{.���8�I�E;��I�9�Lu��~��rALdg����e�o���ز��5�zA������m8򤦵$���OC2E�76EB����Rv�]]y�����jxs���z�y�i�mq�~3иrI�H�=�c��as[��;5ԅ�ޠ$%�n
��3�e�nS}��t���hb����r�]�?�`���v�S2Vu��� ���ūE���������~[�ԣD7�aUF�������L(�) ɼ;:�t�*�-gCx��ˁ����6�'NH�Q�� ��@��ly���k��!#�A�MM6���]}�o��jU"�T���ߍrÏdW��H�׈~ ��i�tAAW����)����e�'�`wk��!������p ������B��%���=�3�_c]V��V�������y
�TS�|v��6�LG�rXlxVHYEB    fa00    1880տ�s����?ʲ�t���t��)��2�jN��2�&B3$aO�G�ac��,=�u�7_34�?^��*��2���;��r&���I�FZ��G`
�H<ܚu�B9�^\9u$J��C$���|�f��'U�ɵ����ও�Z'Y�!��ze��n����}b��S�xp�8-�ɚ�˷���GI+��$Qf�px"�>0�+ՓL�Q�I^Zb.�e�<��}�I
��Wm�K��8]���H�'6�T��G��9� �����Ew2�o_'�L�j�_���)Ei
l�(�u�r����Oy�T��U�m0�(k��U����E�#��@@��|�^\Ь2 2�p��;G�b���EW�e2Y�s�p��|�q�ؿ��ch*KyGo�8O�T���U)-�.k����%�;gyc�f��N_�v�Ω�m�ٵ:�@����c
��#,�f=�Ut9'*'������3�!�~R>�<t%�/�r���ö4S��QY$���n�h��R�o(I�8��q�^2	`~�����:1��;Q`��`p�%3>���ƀ�Zv�������U��֤�Mm�Xx]{�Xm6sD=�^6�oU���Ց�/&��C`��M��#y�˞�k��-V`h(D<O4�78��.r�I��D����s�߾C��;�p�I���gn)� U��4*7�а����"V��O�a���d��f��)?8w�__�y]˹J�MQ�����r��F�Kƴ���V��9L�|��R8�r���A�UB�2^;eP���?4�Ҷc��nEIi��Q�����b4����7�UJ�D�F!Ԙ���]�|<����B��m���zb%PU8R¡I�$�uZ�nҴ��A+_C�Tɇ�+<� E��6�(l�Ϲ�e��S#A���SÛ�: ?mi����ū�-�¹k�
�T��@����!`8�Y��P#v9�?u�U����g�tD�_�z+�s�_�5e�0"`t|���C	p$��{y?}Ώ��)�/�]������bD��@3R���>}�{�(Chz��9#BP�/�����+3MuX�Ձ�[�΂�D`hu� V��I�R7W�:������i�����3�Ev�0��zj!w-7��gK<V
ےr�S�7�*����	��W�A�Y�_5�u������R�:O
��&9}S��&fu+�@�cG��2��iP����t���Bx�SGI�I7 ?�b-n�d\��ZBe,E��� Z�e�{-ޖٵ����y�4)T�7c�fg����Lz�~��I���>�� Xp��&�"�m�ja�R�~�H�xȄOl���i�-֦�n�;M�z_�R�i͟Њ�˳�琰����ׇE${�%K�H�dʝ"��g�.ȗw"��s�z�8���Ƃ�z��	s�^f�XŵM��|��K���=���������ci��=Q7}����K
�e�XB�K���mt8�4wAVI_�X��l��|�k��lXԣ�f����1����ޕS�_@F�(um�ts �[_����u���N1h>���q�x���c[n�nQ��w�#��ºj��T1R�e��䅮��l�R"vn�JE�6�̥��ė=��b�[R>��E�n�E>mАq�����p6�Z]~�����t
':(Wy�FB�y,�)bAT��E�sɍ_��&g5h�X���בsb;�H��أ{Lb�P���n�?ƭ��[8=��K:�8Sq˖2�.�9"v����"'�%ۻr���(�Š$X��d]�V�Ul�a�	���p�`#�ͤ�'�bxdγ�};���z+����D�����yu}�%""�۱��~I��lB4eu�Ԣ�����c�|��M���#|3���
n)p4M�9z�w�	���.[	,MX�e���I?3��K� �����45.�Oh$��A���S�^z�k�Ɂ ����&�(��0N2��Z=�L��SP2�NO���~��uP�����롨$�n�ջn.��"N���u�U��J7���A���J1B��	�d?G�M�E|�Ш��U$�@�.֞i��k�J<;h%�
�x�::��S^�>�9�pʦ�'��s��d�H�Ŷ�hq��ki�!+�^��RR�E?A������<�(���v�j����G�߭>��se�E�h��ͥ8e��|�h8rT�** E'Φ^�=���X۰t�iUH캧��K=�?W�{?��\�P8�|1���L���f�I��L�XA�&$��A_C�n#}���N%��0�����JC�|�:�ᦰp�����qING�aã� U���_�u��z"���K�;��$��F\}=V�
�9º2��b��2��ǹ��i4��g�J��^Ր�]�-�"WоE�mhn�=�9[ۏ�(�o�|$�B�W��~p�8���듆3��0���K���Z��1{�T(��{5.cz%mV��Ӑ"n�YP���F��@�1V�rOG*v�jٺ�[�<���������&8s�<�mވ��F���+�����ǉ=����;��aЯ��kV6£{K�e3(S^p??:��+����쇛�,��l�zo�G�.���K&���{@IG=tX��ck�!�I[�=YH?  3?$���{t��������3r�������Y�kUd�� �-EY�,=r��S�����[wS��^ڌZ��"2���o����$/Ж�������!0��P�p�U��(>�G�"8��X�]�k��P+}㹘k��Z��Bꔂ`#N�3׺���v� D��|	��c���yc�\��^Zn
�c�G�M��Ѭ���/�<�d��"6e���=�����+��o�~�KǳF˶�w�D���@�5�
�
JfK�wε-T�O�������ܪ�"iv�%�E!��i_���5������{_�û�-�-"^�>W� "r����# 2S�r+�\˦�u7:�>	��Wm��l�e��<7o}��Bj�M1�-�D)��Үlb?�k�u�j�|�SPe����)��B�/�қ�^��y�˳���d�ǽ>��	�~P�J���d�����\��g���P�U��]�/=>͋�'No<Z:�i:�A�/�4
zD??J
N���㾾�zc�\^+靇#t6l��5��U����Kq���?���jbPV����e��?(+��J<Ob����q��B���������,^�*,b��B����PC���K��� `�2�\�5��v�A�LtG޾42J���b^h����U:z��ٲ�V��ɔ����e�����n;��_����m-���2��aZ���S�[m4��"qR�����	C)wS�(
����
�QӬ*:��$������@�iu*)5w>x%�"J��=���c`��b����?j���u$i���n��Guq4Q����r���X.�bß� ��%{J������P.X:D����kYh�n��;�9���"d,���}�[�4�]	�֜K���
S�W��&�̪U[l/�$v-O�[�kK;��٣�4�w��{�,ĵ�L �����y*u�mx/�9�r�31
ȼ �����}�?�ѧ���E�/���y�zx�*�+�H'kWvfS&�v�p�б`W�Sx���!n~GS8	S���y2�Х�ݎ��Ft���M�	D��H�_)`V�xx���Y{a6	w���S1�>r��#�." �9_�)N�H���8��ã�P��0�����kU*���3#�L��3�۹q�jec.1�[d����B+>h��ye)5=��[�jD���lT߫e�+�J�Ȉp����&b$�[;�~$��"O_R�P"����g.���Ik*;�ʚ����4�	�f�Yl�фG֒�*s����c�n �i;q�8�3��e��h�`�pt�S)<�gԶ�
{�:��b�x�lTd�u��{��+��o��Esd�ϻ�"��6-Tf /��ѝ���T�uZL�i��2�����SRFU�g���Нϱ��k,��ˈ��C�n;�5N�bfT�_�~#W���b'�?0�I_'�����]��1?�QZ=��֪Ě���Ka����4���^�|�N}i����s.r����gt��_�������Ȝ���4�<�]��n;Lbܼsj+��j`��.W��(J:��5���gy�,�M�7F��1��÷6}�2|C�ź)hD� )�:��V��3�d#�˦�m�D��#>�5��8��p�f��]�F7t�(^�����8��`HZ���G����\0*q��h?q#g���ch�D�ؖ�8�g��E�;-�S��.���m4�nz�)ڢR�����m;<�;��d��W@�Wb�i��[��؇ŵ�zF��Qˉ�2�y<XO���tL�P��2��;}�6��ʼ��~o
��~��t����{���B�G2�>d|!v���d�3�HCl''��J�I�+�>z>ܸ�����o���
��ъs5���K��]�l�U)�����[0t]�f�0�t��t�/�B0�|�0��gd��� ���˄�%��������=e�#`��ȫb�)�-� TXOй�(��ÃF�e�(tw��W��$$c�n7����r��o�)6}��W*@l���=�w��QOs�1�n�T��C�8�`��%�PMhܐ�h�3~��f��r���2+:����#%����NϏ���N��z�T�b��Ez��rHT�����)4�8�%�-��:��	G��p�ߴ��qo��r�ch���C��ZC�a���+~ܗ��Q���
P.;͖���YD?{�7r�#�vv��:(,u�ϸ!���p[� e�nA�O��q���V���v[���C���:�I�m?X�m��lnD0sI�b=P�8�'���I`ٳH�7��>�܆���4��6-��+����O~�Ww�TڲJL����u�-AB�2�,��4��~�W�W��Ǎ�*>�"ڃs��;�tK�,�jU�X�����\Ν�eA���̾�Q���>k+6�E1�Ʊ���[qGȅE������j2G�D�&T�(Pg��I�Ъ.%��a_w��ZV�W������BJ�Ϟ��a9�8�j�8��;�wo��nF�5��ND��Xo7����3��
�7�2|VNu񕸮����Bӿ�u�������i�f���^*�*7��%��-���u�S��f~Q�� 0,�Rsf-
���~��[�$	�����V������ɤɬ�h��^��·y5�ZW�o���0@h.[V��1'N�L�
��\�f�\��R�b�L���_FHm>i���@K��t�/��0o��@>��)�����a0*>������N$�yEY=�bR�4G_Q@�'��+����6�D�i�N�T�4c�j�{�wQ�KK�#ӳ�,y�����,b�Ycq 7U��=;Y A|�3RtcU��׷���C(cm�R�1"o���S��_�(N��V?nī�!{�ܔ�}&gR�>ۻ�0 =}.���W[�'�Sj��1} 	np*�bo@�b�ɗ>��g�<0�v!G���r W��n���0{w������{<n�R�"��?Au�V���,e��Lf��-Ǎ��8.�K*ژչ�Z�� uESߢ�o�4	�Vg!-�0���7�Y���U-p�0��gF�ob'g��³"�#�@��N�2��\I�H�2-�su婟�
�C�z�
9�ɏ�a�#�����ӷr���(δ�4��]Ay8f(�����R���0���Dk7���G�nE�T���𑗺U7H!(�dX���x^m��4�	�4%e{��iv!�®�g@֡���M� N�Bd~�1	�h�~?
�!�jTwR b`���fɸH֥o�[�dܰ��fG�ZC�/�Ps�Vkv�g�hh��]���[�POc�����"�;OlsI܇"
�k�� ^@�S9`�����Iso�X�q��s3O
�]��Y9�S�b�,��c������v�Q���;q�l��G�1v[��~�e%� �ԕ����Sh�@P겅��g>+���*��:Q(;W����侧g���W-륗(V�1ct�.��	_#]ȸ�Q�����ZR��`���E��&�O0���hm����a�ro�4v<T�����y2$�im>�����~�sա!-��tc m��~$��M=f1�B��1 �7K� �ƇU�ιi�-�Yަ�y�>Hw�� �cz婾����o��Hj`����/xXlxVHYEB    fa00    1910	��#v�IͿ���~�.���暫�/�<�{�-��7,$NwS�]��M�Ո� \5�D�g&s��_�tr��m�ʵl)�QF���_�fƱ��� ��X�6����Gw닥������	6ヾ�qP�B�h���g��Ѧ��"����za�\���ҵ������ 2}�A�͍is���4mA\��a�u��#�SS^o�oH{ܠ��>uբ��'#�X#��D�_L�)G�'����{��"�ְ�nѵ�?&�U�|6M��N$
)���6S�vܷs{H�a8)�|�w�o���,wwۉ��E�����U=7��!*�r2?�ք�4�xx"���朐��� �<4�h���<8����6���w�J����4��ǎ��� �!s�cu{$�)x%��)��~q8����������{.�ۙ��S�>}�lrsssv�g��J1W��A��jc�v���o���r��i�ۘ4���E�9�D� ���l�h���>��궶A3
ƷȺ��~�b�X_���sJb��� �%�����J��u��(����8����`�蛒����Q��t��v���*1�́\�O���`n|n��"a�	�4�8k�n�A�Ƹ��mү�x����%o���<��w�!Y]	���vnè��V+�S�E���'�(D�L�	��y�.Xdj����<0�]pd�ͳ���Yd}f�F#�a1ؓ�u:��)_�������T��-�HjӾ�I��
���������ʱ�T{�ID���^ݕ/ܭӫ�Ԁ����>�;ed]S����6Z+��F��Z����6	;q��0X,�QW��֤C��L�	���:���Lh�����A��h̻�y�<G]U��T��`OIz��a̔�'��s�|�H<��?��E#w�ͤ'w��Xf���.%eN�ә��C�-0V��5B	H�e}�eF��|�L~n}�n��;��ݱ\9V���<�:I�S��!��L&�<Ț�::y�j��4l��%m�QXQ2���_���S<���X���[w��ҪM�hS��1edz��ǽ��l�u�I޻p���F�^�}<%�I��ҩ��L_[����-ƛ�;�~)����ĕ=%�������P�|�܊�o Z��U��H�����}x㠴+�
ԫ?�O��T.U��s~���h���P�t۫M[72�p �8����������+�QӠ�B�gB�E@[�D0�#@��J�e"w&�\�?�C���1	
��R(w��.�wh��2�Q!��
h�P ��7�%c�*m��B]��6>כ���v���Pl����L����^��D������ʷ���͵è��6�J�Ήe��H�
�7Þ]�f�uQ��,׮�i�3=�Zm[��[�IߵM� �D�B� =xm�!L�S��������%�eh�`���^U`1���Wg����Y���R��(���.��T!�h��k��f95�8�ټ��˚�
�B�.�h��7����<�R��k����V-���EM0���ꊡ��⌂�w�A2�V���nU��RF_��P�]�p؟�j���`Xqj3B�rexq�&kț���X�))�<�U�����Z�=(�-f6��iO����i�V/
��jg�\�f`1Xt�y��S���Oά7|�����{X�q�	����q���!C+<l[7�>TI�Oh�ױ��l��b�Q��L��`2Ob��v��L+�W�%�Y=u�H?���éi}CŰ#i�h�v"��p�8֣T%�$2�����5�,i�u����@�gٿ���\E�� wT:��G�������DJ%��o�B g�� ���fיQ|uB��3��<�~�u�SN")՚Q��Sg$u`9�~��N Nv�xuJ=��de�!- �Y]D��\���z�I@.?�E�+g?5p1���c��6l���ݟ)i5q��ơ?���i�Յ:����KT�,�ʤS��z��4Ю���p�^Z��'/�w?�#�Y�{��Q`�0~��uf(6�4�8�9Is-�=l�Pg����̒�����Qc}q�sd��b,�!�K���}���A=�����vX"P�n4H�x%�Y&��V��n�h�(�b-QmH`%xE���<9bC1B��.��S���rT@{Y�7�1�}k'�G ;t4]�7s��:a�t��;{�\�T��}�a#-)�~b�&|���`�)��q9͒��'6"&gᣣ��~'��k�h��%k�o1D��ڬ;��������<yO;�J�������KKQ�V���� �HN_[�o�s{�y��� �4�G>б�M5�I�R��e�[c*�7Q�`�8(W|���k�����r���0��^Z\�%ϥ�;'�	P��LJ�!	��Hl�)� �d+��x���Jz���+�ҒE.��m��R>�>:�xM���	���k�'z���-�OM�Ժ"�KUc[!�P�y�,�V�N����5�.�E8�P��D7~f6(�/ )�\ߵ������Sx���a�c�BtZ�sD����E�$_"f*SB>Yf�V::+:�����`!�3��;��$���pps����yK� �`D�J3����aT��6E��Q�2���e�y�Q�4ڢ�"Κ*��.����C�����"E�mV��U-��$��K��R进�Q������Y"č�/-_A�(�SQ�`7t�垟�EkSն�*њ�HwT��^ (��m�ͱT�����Q��ew�rC2ȵ��C�tǡ�\p�<eq�7x��E�r�0��;N���sd��6�����Bd�R�T�}��Ƌ�"��W�^�̏��睄�G0 ��[�����v�IΫz�٤Ԕ-g��a�7m�Q�(��ѱ�b�1���CC�0`�;d��hNc��}$V0}ۘf�Ҋ�����h��=q�w��p�1/6ON~�ڭ��S٠�'�Ѻw���D�.q�\*#V��I�&�X	D�M��XӐ�\H�����#�
L���_�MugNwi��`k��me�����-�������7�JeCܫr�,Ԝ\Q���@:�}����һp����������nqA�
T�'�$y�p1*�|3��iFN�1N�`��ID[�SJ��[,,'�~Y@2R��/Q�p�Zy(Y���8o�`|4�q"ς=���U�#_w`=��|����ع(<��B��8�[8e��mLiNϲ��i$!v��̯dɕ����B�� %�LSVg�^��o������M��*f	�����4�2�|cc�ψM����`,#�3?�&n!��}%ϒ�v?������0�.�@SNt���`'��h)�w���}!�۴����ʇ}dAHN�i�j�W�{������� �G"�b�R��$�����˿Aް�A����2P�n1��<&T����0w�� �i4 f����z�aa�h�!�P�x�Jy,�j4��$���K�x&�m\�G䷘�ц�P���y�j�(a*�(�^��ɧ��gO� �#�#q��������_ZB��S��ۏ��7�alnR�m��ȾrJt��$��������b�.��L��+�)�.�\�Af����YKU!-}�%؟���%�AL����%kFM'@�j���Gm�78F�ݰ�ɒ�U/Oo��ۖ�M4#!�/��gC�J���)��[�K���J���U�K[�b�J��6��=�����"�1��"�ħV���&O֙3����i8Nv�4�Eg��Z�|��3R�K��"w* f~�<�:9p@��1��m�}i4l��@�=��Gt=Ad��ܪ=;@'	݀�C��p�v㶌W��]��޻<q��ԫ��F(��1�t���?���d���%��!61\\a�`+<�yY��_|0�nE�w�)����FyB���ۏ�ԋ��g%4���r� �~�ɑ(@�V���#�>Z�u^|�f�)>M*�v��%��l7i��zv�B��kF8�������wH*��
�ĚQ�`�K ��bn4f`�Ѽm�����b���.�<+[|��4� ÷]i���� ֈ�u�ၙ��� �<�4�&�Z	Z;Z:E���1���2�˔�:�zͥ�u;*��^�U���5S�fJP
���b�H��u�
����ƽ>�@g�^���l'���#]W@�Kw���wf�62�3��~���$J����C/�\gE��i��U4��LŠ��ڎ�-�5�_��A�fP�[[|��v������X�|t�K�sM/�x�Ճ-�͚��.�l�x�#�dpwY7�= }=)�����L����-}�T�jsep��^�:�h�'"ٻ#�>�6��~��øv�wK�a�r�g����dh��K�b�}T����R�f���5|/鮉�Fh�h?z�~n̿���O��9ìO&:�Ϫ�vq��k����s����2��\a����������?4W�T�/Dj�-(���t�+aR�����e�#�����J�Ki%�k��25���Lֻ�.*�fj)�H\�)R�	�eS���<#���#J��G\�5�r�@ߵ���� }NoH3�7ۉ��A5���@*O��O�h�6\��l���v���˘׀ ��l��c甁n����a	8I�|+&�-0�����_r,��������a����V6d��dB?lHm����k�|�qh���6���h�����/�I	�Ȥɖ�⠢_�����O��*T�^\�w�����TӠ����  �W3�ؓ�e�j��] �y�ק�L	 ���,h�0]�_0��`�+������o>�O�&Be��uG����=����^�.v�(�b�$u��Ւ�&�����G$�3[+�t�j��P������*,/�@�U�� �KT�ZA3֦���pMVnl.t[�a�����V��eM�1^t�\c1�
���$��}:ϋ�}ԉ@G
�#:S!/k�gu�|\<���$��g_�e>S@�I|K�����.�B?ؑ)�J8�G���佸�&'%�9I>e�����oi;Go��:H�֭
x@KK�n�ɘ�|=Z�{tl
���64�g̍6g${�0��s4^{4C�Ӊ�����
�U"<[��1 �P[nԇъT] ��KpOK~����%l� ��n���ObS9�&����������PL�����l��1�rG[m��rЀg@�Z�s���l�R���Z��	���:��JTө�b�`�
�m
ܣᷖ�1oF��C�<�*QT��\�N2��GM�d�)k�db��R~���������:��W��1�O�i�$>Ϯ�̞� H�ک[�j�8�4s�7��}b:%����,�*�^}�/ꈾ�\�_�o̽e�xW��u��E��5$/wC�)^�)����X_MmI/�����5m/�����#���.�������V�o#�s���5�a	�Ӆ�y�&���5�q���$*:�Y���R����c���756P�x��~<bOL���*��L����P�BQ���݆)N�>pg���Z���N@2���"ڏ��r�3����㗠�(Lp8�	o������:��?=/���Vox�7�DD��`�����\ŹU46��Z�'o��� ���("ѳ�F�a:%�A���kZ�����]�ߐ��L��j�[M�R6�������\詿�I$����p��%v\{�s캼/=g��|�X�j��
�*�����|d��)��R)VB�P2�����/RbQ�c>�����6�_��'"d||CFW��G�b썛�qQ=e���<�TAf:X�A�y���Y��o8� =��N�Gs7�̪�d��d��
a˜������hF�4M���������T�9#?� ��/sV촡������R�I�-*�+mów8�u}r�Y��[���̳}�k4�Wv�^��2V��>x�֪w�3ߡn�	����S��>Y� $�`��+����U~�Ͱ�(�ʎz��	�!��;�5�?+�����z��?(�.�c�[ւձ��x	�1����/䪫j&$�"k��;N��y�{��үJ�A�Nڠ�	I�p)�H��lϦ���]�ä4���9('�.^Қ����~�ź� $6|?쎷F
<S=Y�%i7��iU}�\���9j����!�
J�L�����R�J��J:��ј�!���.���yS��`��5�*��js��:���m�# '��.���>$34A܂�5S_���L�g=��0�8&l�Hδ*O��u�Z=�U��D�L�c�VP�`�x�o雯��O4�ၜ?~)@����ע�'���ז�6fXlxVHYEB    fa00    10e09UL�P�m����3F���A��w����eo�s-����>�?�+EK3�e{=ޙN*՜�1�U���D)�m`,�*2�-�L&�X0W;�����f����w����&A�P���c;$����M�Z���(�ҚA0a�l�{n�1ӥ�<?M4ĢE��m␻U��6\�JczI���k��U��13�* 2Lx�|�X3�6�!B8fTM�5�>����+�LO�:\��#��ۙbi��U��٪U��Y�th��a�x&-�jM�1���BJ�(�R[r��"u/��!c��줵KǼ!�<$dj�~Bb��VV���!0�׌���6b?�����Fϼ�\�����;4�&eo@���8�1���l-��4�<(���,�C���*D��SS��J��y�)����o6�lk��=r>��Â��Z�|Xȥ�U�?�2�.�}�4���;�:j|T;�[�Q!�i�lmc3ئ廩�
����J�7�O�:�u}և~U-r������G�A�] ��Q�U,D3�^��IYީ@��C7�#���G-�m��I��q<�M�a��W��`�_d/���7a�w�Wwa���ވ"p��t�[K>X=� a)'���Ipp�-<��=�����.�{X�0�L��<ϕ]�(/k�A��c��4#D�=����)��� K0ZX�ս
\����[�>-���1<�?�g:���@Bw"�e"e�?Ԡ�$�a(jg���r���Ͽ/����%����L�Y0��Pb�$Ձ[skYG#��������)wJ"�@��.߻qV��.ܳ��v��NK䵮M��t�_�ӿ�%�d�lE"��=a�*�?��F���+��MZ8�ا�>6�f���I�OѶuZ�xY��QI£G&�!ä:�F�rK����;��R���	K�t2���ݐ�y�=��V��>��z���/IEXbNxH���\/��Kj|t����Q:���|@^w|�H@s�(v�k��k>T�s/#�����u6u��9 �*�v��a��>}X� pM���l|����=t6����?�9�y��X9|�%�gyo]�̾捘א'���Ei/]��C���K��G��=Ǘe�R����n��f�_@M�[O�5��AE��ɸ����T!��	���Cy���t=5]��W���LG�D����[���qfJ˵�a��?ʴ"����f_ ~a�1�"�93����
C#��Rd��'� ���±�5�p}�<d<�!�����V��76B�Pv���-���;;�����@ߌ�"͡����r]��g
R����@�̶��2l��eb%�W��L��w>���P^w�C��wl�a������%�-G��>���a���R�F4�w~�#��1���W	�l����&�ӨM�ܞ�7*W��S�`<��m��ɓ ��Ut�š���T0"�;d��7��[�!w�PBP�>,0V�tj=^��g)��C����+
��ɝ�������^nWh�D���U�C%f%��vlQo�>�*e�:�@N>]Uq��������ɐ�jMF�V��}��2id��f�/W8�4�cP��
���6x3��(�t�R���!I��ȑ#����W�"��B\H�b��X˽��Zi]'���8}Lq��R�5b��>mAM�Օ����bO�M��>�y�o_e[�BB�qWʴ���5������Xz�Ɓ��d�U�\eB~BK115Ș]�$���h���.��RĴ�>\}ON����:��R��wH�}}vņU!Sf�`��}����#Tv~����b�B�d2'%�3�JL��MI�a��+��6���FqOy#�LKO��]�Em���	�S�ŵ$�L�b�������̟��&w���]� t���;�3y9���a��PW�|
�zr�n����Z�+�N4'w�0L�l<�,m�/�(R�<�Զ�uʮ'>�*�pr���=��.���]�t��1�7u��:=�+m�*8������󮡟|���Li���>�s��L���"&qz�����H�6�M8ka�x�}�S�1����.i�� B���/����ǯkN�?|oE?{�Q��r��.n<qc�RlX<�LK�ʭ�Q׭2EhE�-��B����D���9S4�	�"�Sz���Ѝ���̴ä����1В��PX�����b;E��.7'V
���c�i��.�q��/�T��1�0�� �p ��qo^�z}X��QjP��������=�ߝ�Dٯ���������Q����8�:��sUpC�:ٵ�v����#W 6�m$i5�4������
Q���Z�h��_GO�~@�X�g�'���V$O��6������{��W|�f���	Y�������l.������M��K���Ŭ���q:�d�@kY���2L��{��p̂��yh_z`�C��;n�SJl4 G}�k�qxvs�Ƹt�ZU���eݥ������0�RV�0ov�t*���K\_}$�s�?�ݖ�l#�4K�F�E�'�l�kFoV���4S*��ʦ�c8k�Hć�`jX^�z�w�+��Cr3p��1��1��q�YU��"Õ=K�
pQH�wK�$^m�]��j�x��FS���z��h$��XV�0uGv��[B�MӇ��8��Bj���{"���$���n��t$���$���N��
>�S˔�Σ��"��M��W,���P�k		ƀH��#8�	������o�r�J#�%�ʟ{��0�T���.����&���h�4��,���1�2��Ԓ���*'�Y�~,o��H�%r�D���K�ǹ��g������f��|Ua� Z~�^�+�0i��!K6�6;u�����u�
X��4v���z5�����$�b���i�f�Q�%�l1���m����9�#�"|�s���C?�_Ϩ���������`;&g�s�iY���������4Yn���D���#��x.�mR��e�a� �����/���'9y�D���ky�ˮ`�W�Krf[:&컋a=�F�\/>�plJ����f�ܢrE%����B�{!T:LV��]�z�Ϗr�,��ޛ ��˳w�'M�UY��L��ѥ�,3����;��\S�=�_5p�>��.~�GS?R��s`VQ�I�@ZϺif
}c�U��zd�V�C��?�m����a��X���1AȢ�XĞ^�[���B���*1�����������7>zX�tL@�J��=>;˪a6�����8{��z�?UW���.���Xց5q�T��j�����G�Jhך��O��-8wc'�ސ��n����	�׿�9�U�Bu�̠��[K#M�0 0�k��?8w�3�h�$��6�����ZW���?[���S�[_��3���֤,y�!`v���0��E���X��Ո����w4�<B^|���{E�
z�!4Ttq��$@�{��nx�J���RL�C��xu-N �j�
1Qx��8"�/^�ʕ��e��Iӻv�?N�8�%E�R��~�X$�T��.;���v5_���A�͞�%�q���4Sʴx����
yP�kUiC8�ԃ�5����P�����̋wɁ�P�1�6%؟��w�쿛�j�,;�
2��� @��Ï>��_%�I���	.�|7
\�}��3�GhNTY��,i_dX���:\�<�qR��	��J��kKg�@���?��dY��( ��ZP!�sI{����Zi��9�Z��r)�R<3�<��SU7@q�ܥݗD(ֆ��K��ܮts��3����!��D���[�z9�{��]�!�E�=�c�UP$U�w6��i�:�8�����rj��۸�JM�v�N5�]�����)$?'����Vt��
�2'5���Mk������5D[���;X�&�v��aH���!q����/OyQv���@6~�ߞ����H	�5�q��.J����;�с7o2��@�\�i,̳�F�]�v�$$D[��i�@82.��S�Τ}w>�A*]Csa��\�	��|!�A�5	��ז��|ɀ���HjsI�w8�@�T�=��{�9r"�vN5��v�4���m(L��:��c�<�9A�|�W7�LPa��C�D}�2�V �R@<4M�m~~u��c��RJӼ�۬,�M�ظ��Y_��y��󽥎Sh�u�h�t� ��E[3�����ԭ� rY�en��#%�8�]�.z9D$RWq#�A�E�|���{���%{I��k��Ԟ+��)�|l�E���k��'��Ќ�I$�瀣�E�[M��t�9F��k��5g�!k�TU�)XlxVHYEB    fa00    1860X�eغO���8��Z�	ާ��u����z1u�wל��M[kG�5~So{�X���%����)��7�B�E	<O���H�%
��y�^6@q� ;TZ\ų�-Qw2 &uǾz���T�|�1.�{,'�5?���	|��/+�&\h��~r�}��9������c!sAB�H,|L�_a�:��pU��tr(�Ƒ���
S�o�H�
xx�ѽ�(�a0�j�������`�?��Rk����l`S�H��~7����P�A0L�S�������}ь��uDR��33
��z�dC#��v��U�L�0��,ކ�P�������	=Ӈz����`�n}{D�'��Y�B���=�}e�M���O��]��c�G��0E^�
�p������^��瞺��NÛ}Gz���?v��9�%�/F��f#5W�8�i#����A?�z��*%R��Y��/��"+Q��I��q�\u^��b�����&�����t��q����w�7*��WF���i�Z��O�X0qJ��Ov���^g�$�j4i<�»$���b}1VHZOR˿�(r���C�y�rW�>�ۺ�%m�_��FP ����{w��(�J�x����\��>����đ@��&TuV���]�R�S�$�ޛ�{l [g#5�T�?�*�E�����H�ҕT(Y*�xȦ�rX��h�ӥGk`3�������`1n�2i6����ze��NL)�ʋ����O�Dz�I
����Lh�5��ы�1�i�H>�5�O��}J}��,�"����\��.i*O�� �,o�6���i�(�塧tż��\(�=b,�@��r�����V�T�/F�H��i��Enɵ�Ct舦��sY;V�q���։V�n}�ӏ���&��YRM`$�(s�>Z��v�cݒ$�,w+�(-���w�Od�^.g��ŝ*c��t�`J+	�NR�.9g����i�>8���.J�.�1AID|��ϰ"��yQs:�A>a�L��Y��AȝX}Յd �Z\J�O<ZE�!ڡ�ztks@�4��[(,�Z�`����(����{t� ~�ܐ�A�E�'�.b[_KD�Kݜ#���f?���[&�b�5I%g'�Ǐ$.ҭtH�b!��b������D�xY�=x���o�NP{"��Iک_=���4�Q�["��D�~�.�/��t�
�\RjdȦ�qW�b�պuI�@�?&����>G{�h�����{d�w�����P\O�bx�O�6�Y�3�?�����Me)[`�:�M���1A@�"�n,99҉(D�L�ͦ���VF�N�]u�&�*�M��@�`)[m�bQg_FD�>�;�2,��{�A��v�>��{��l���
�8��sd�X'�}��O��t�aoP~����nZY�vr̻�
$/��j ��'	FQKd��
�*�/�6qӿ$Ø����x��U^���4�{Fkjwj{�Х�Y���Y�[�/VUC��+r�&��E(F�s�g*��M�\�@��5@gՌj���*Q 9�]F�r�P���Jɚ3����cN�ݓӄ��<��R�>�l��(���Iw��3����
��S���@3c�ۜ�����Xy�f�l�09<.�`tv���p�u�P.շokā/�}�`��g+8� �qsl�;`M h|���Z/�=����`m�<O��*c
�@�%��#�o�3��l���B�Fy�q����k'�%;^Q�
���^Fl��-e-���Ւ��7f�H�n{�)�xn:X�����[0��5��󰪾��>�[���*���Iw�	�2���C�3��s�Q�8߲;���!?*$0�'ղ> Ʈ���a
I�[p�)s�����Ru��!�\�Ͽ}�������}r�M6�������Je*�^���`��Jh�D��Smc(i�դ$�=
��P)�+t�5��C��T�Z/:�y^�~�%�du��Q�s����s.n�h�f�PkϬ�ᮞ�Z�6Qh?�]"���Ԙ��J�T&"/�fH'k e�?cɬG^F���r�eawv�a
���!V<!A����L-�Qdw��\��U�~d�
zG�=��T�m:	��+�� Z���P�\��>b����I����J�%	��Fd���G�֧������"|�;�����Y��	��)�*2E1k�㝿{Z�[r����5	�yۦ��B<ݔV`@�m:�²��h��b!��_���P�<� �������Iئ1=r�o��}<�hb~�L��O���3�d]��y�\@7ꤐ}G�eq��b8)�h�S�}`fgf��1_�	�Ȧ�����n�y,O
 �N��͚�^�c��
�w_r��a��;I`1*^�GM�D�4�cF����&��T���A��pꣁ�݈�Sƙ�v�����9�q":��8������9����92�p@@�eE�rY�`p/Y#R�x浱ުݘ�E�D�0i��yq�7����z��C�r^o��ma�c��`��b&�)u�{�t=�L��M�&����j%bH#�i�X^��kK!y@��	Fr�ێ@�a0�H�)���b�	$�3Yܬ~>�h�1��W��8�Mo�Ӥ�r�,����I'�ie�7��]J(����74��W�Q��8NȮ����x3T��NXDSϩ��5*� ���t��Y`3U��[[�R7��|�TK)��K]�N'!����qLk4BkfJ��9=OM؂�CI�5������	��� �������QC���z	��:?*ӭ��#έE�Z�SP�q��]�M�,ǆ����-X�8oȒc�;�Q�u�7��!.�B�ic���-~8T
E1U+3���I���UwߎG�"��,�S�y��xo��?�Tqm���?^)�x{[]��tc��r�[��)KgÁ��&�0p&H!�gw������)�f��`!�VIG'����bn��������Xճ�>uo�!�D���<�	{$��H��^F��KpcN�׼~�bg^�Jt=M�Gɚ����L��B��$�XXb�?��gF�7�؛Vg��(���!�M����8r�EG�*-)�"dk�nV�rBU�%%PD33�n���wz&u+v��>G�[�[�d����<�"�O�R�1��N��	������vp�vGq)�����)<z�+J���<oqZhA��CW����������� �p��҉ꓑ�L��V[�H��q1�Xܬ�{�4�x��s�R��{k;�1��4z����Sf�Ah�܊�|�/��	b�D5�s2r[�5�
��������1����Y���;ፚ4�h��x����ê {Gl���2P%w�}t�X�x������	�wE3ױyW~8�c���d�+���8��4a�fj���6R^��fF�0e����8��
Jt��h��m��3El�Z���<�&a��"9g.��Ю��o�=/{�F��^]gRԟ2�q�3吨�\+c��|	�˲5�^_jpb|B3��>$ծ��N��o���0d�Ȣ��\����4�)Wͨ�G���R���"'�����!a�a�P]t]Y ׂf�ʳ��A��^�G�odw���q�`n9��*~Yna�C
C@�%Ӯ��h�69
�Yr���6���K���V��#��[Z؅~���j�F7¹�C��Fh���a(O��E��%xbT?@m/�@�ҝy���xư��ƒ�6����{����F�ɯ:�3%��@q�����M�D�n�:�T���q�<5���:,E���$$� d�#'����+?�h�����f[tR:V<�摡kS$��L�Jۛ���7S���8eS�Ν#9�����S�`�=�Uw��E�d��?�b�X=ӛ�&��'%����
$��𾖿/Nj;� R�"�ќf��ODMVE��^��r\��!'R�ٵ�F��iגv�b��P�=��qn4����e!=Mnǂ}��3�n��
|�G�WK)��|s$q�2v���e�^�����8��[OS� ��au�M�(�E�!�n��	�v&aS�O�F�>t�M������gw��C�����ʝ�O������J=G��ƬV3���=�(2lI4�)��;��|.���:�ELus����6�2��QB�d=�X����>���6p����3�/��{�\	��/�6��L����$s�I��].�-�5�^ 8��$M2W��ف���h��s��j>G��`H��?�Y��`P�E71"��p�%�!a�u&��u4���Da��a��t��(6g�ڭC\/KfH�]G�υzAd��Nr6P� ����|ա�)%���A�W�����t���'nJ����9�<=�P3S)�ƌ�>��	��X�;��~6��f [��k�8�-0����s��7����f�7����S���Qxm���f�C�d��5h ����~��0��s��ӎ�5yc4cS]�3��]2�NJк`�x[�?^��4.�1a���̆�t�?�u���&����ԋ�8L�b�����<)�!	�JX���!&��L��>2���eZ�p����!q�L�ˋ����U�,����i �О��p�3�Հ��(��ݥ��{���j�7M�W�py�VD��6�J�43rhn��k5F�0d���a�}Z��z�"��ϏƨG�!/)�U~�A�X�q��Ɛյr��cl~t$��~��/�Y�R�i�K�A��j���酯�Sb�X5Y4Cñ]�B\�'�5fd��ﱙ_��ێ�^^k�����������9boG`M�{��6��+�ջo��R��T��e~�����g�J[
�	����^
��b���s���;V~;��Ҥ��ǅ�<�g���N�RL��GZ+�����>�;����Ы���J
�.��^a\q@1�ӯ��k�IU�%f��p(���I�X�,49.o�e���>P��{�����E�$���!=G/Jĭ@L�.��h�KBE�ͽ��$�O4]����{��rCpv���䙇DO�'=���;����w� �=�<�!#s�+� �q�������;N�H6�]��M�Z*��%E@�)�{���!-�fk��u׊E�Z�%�w�3��!�bzW~��:Q�F%n�HQv`�e�@�P4�	3��ߋ)��#�h?]CE�a��M	�4�laoCw$�7׾\����R����~�<l�=�Jt܄�\��=n��wU���ȗs�`&���έ/QM���Bk���k��yho�������-1Ĭ¡��˭�|��#�3F����Jd����CSv���.! q��6���
����*�Z����b��f�|q��dp��Tu�)_$�6�q����&dXI��($��J
Z���N��G!�.T��y�wg�SYӳ�B�U��Y:������N#3������8�ߠ���~~q�'tHt�,�F`[9�H��->$k���sDT��M�9!Ů��q	�����fr�j��>7�c����8rl����p�W��$+����J�������@3�;�� ��\%2����Q/n_��⪓�f����%��9������TH�i� ����2�r�dLC%�od?[����3Bn?��ж����l:�r��X���ǉ�� yK��c܊4.*d=Ҙ��v��i8Z���/�^A��w���v���^�Рh��Ig9~洵SXNԇ�
?˘u0<����o+@�����+��,�1��Xj	
Z� �w��奘���Q$�h��ϕ�2NYI��z����R���e�$���	�zO�tԞ���o_Cu;���w�O:����Q�uh�=�L9�D(78�wh`��*�C��{X���L}��2W�f��	Y�Bꀹ�q-�P$��6^����}P����������@��+��B�6��҃y779���%x����F
 �ZN��S�"�0��2���!��>'Le�Ѿ(�R��2>݄�(Oj���������%j�� �)O�G���3�h>j9�?i"�������.��?��3�bT4�IH4WBHʹ37"l�7Q�0CS�
�Tp�@��6c�P�����U���D\��-��gC�@�$?�� MR"��a��M����7��m����5�� )�dK�m�Id��dUCD�EC|@$�?����R�g��\�cg�L�a����XlxVHYEB    fa00    1720>�1��E�=;�턦l8n7�_;^�<Ga�j�YQ%��!㺊��>�Y_m����lI�����6�[�9���q���Rp�~���NJ�rȯ����{��	��N��9��5��ytt11>�&_��y���uX����* ��O?�D<[D&x�0&FkNG�,�p���V�/��"8��g�)y��<�O/����� և���xͷ瓱M� ��za��I稒�g��f
|onZ4M�fy	֩��d�]������ +U�8J�dh�j'��^�v�U�E�N9$�Xo�������e�w�뽇�مR��h�d��	4���jd��n����R-���p�<�l}����V�
�1�v� �����2�r~����{��g���#@@ъ���&�$]4��eS���j8���Mtν=�z���A�b���'�n�t�~�;�vSVK�s�����B�:���n�{
��@
E�y�1"���x?G��4��P�(�t��Cr5�1�$�7-D�
m+FČV⎨x�U�5h��݀}7���p3Ҁ�q_#ń��\�E(�G3��A���?B3�����a2��ː'ڑ�⚐5۽}�D����裶���� �w	�����:>�rѱ{�q�ר����!�r�vGT}��LMcX�Ct���7,�t�;���8X��5,uɊ�˅WBz�~4Jϰߕ/����4�-��H�AA��'?~�31ve,Ѧ���	oys1?�U&�f�l!MY_����?Q�����I�]5_F��'�o�,����u%��+�
��c�&<r�/�Y���4�8M�� 2��Mqʌ�<�DP��_��Re^��o��E9�R1#U�hڸH�qԛxս��'����-���:4#�!%%�"|�]��᱒�e�
I�����[5��G�mJ�B�'���&*�'U)��n���ɦH([<3�1���>�^f u�8ho{����rfY&�yctÊR���Cg������Mth�+q�:?v6Tl���K�]ش(��"\^'b�� 7����fB7ngHۤe��pO^� �<-I��X��fwmhX�yD(>�ª��_~����]˪�g�afx�.0\������\�bh��t���Aq��%h�ȃ0]�;e�9�s/�X��HW!�,��ɖ�+�*���s��U � �a�3����븆�&G�7l�;��L��+�tF������w([C���cj���;h ��7f����i٠��K6Ӓ�f<��F��.�V��lS�����mEF�xeX~�AQ77��0Z�xѧI.�P��N���V�#��u�,��!��!�9�m5�]O@ʬd>�G�_�3�<*	�$E��Q�5��!Ǜ��}F����
v��K�2�y�p��|)�����Q`�> ��V�a��H��h�JsP^�It��� �3�sD�U*�zX�f���r�ة?hm��?1Vn)H�d���J��Ȳ�r���_� /�����&��"���{���u�%Q����9���A�a�Jp���~_ֳ�Z9� �"_�s"������ ����1:�f`��Dy�qp�'�7%��%���fs��w�C[�xJ�2|�~��Y��D�Ab�V"{��1��{�bHv�\���uY���
.C	��nҜ�@�b�\h�F�vd->W���t���lgiV�XbT���@,�2j���(O�?����gZT�q�v�'#��B�soc'-���[�,h!�D�x�8�����n0~�}эc�a�-�(�_L�)�CIٛ��M���)w��i�՟��܂�a p{�r��~!-�B✂��S�z��C�i��P|ˤj��uS����W�c��6�?�7`ج��ˇ�_sK�tǎ+s�'y�D�},qO�g���,�ϖ��L�H�'+d��\E�*/��h
��x4|�%���C�UJ�Z�r��ʎ����G�fӊu�\�� ��X�2�@w���b؋A��M���C��t2�	"u��`��f�|�ϵ�����ʚ�����^�Q���:���ԃ�^�ֿi �K����`��X[[�~?㉇�p(h#O_�V�+dʽ8���֪���5�~!
��;!�����%�H������
�0=�7A34m%�^�f�3CL$��M�N�ij%޹m�coT��!ў�鷏F�e$�s�D��v�0��EX�FV��Ɂ~Cl��8��@liK?X�����f�HzG�"�d�SS�K�4�NxR���tA�C����!UY��'��V���ݺM���Pi+�fnJ�2����7޶%>�4�-<%�լ�h�n8Yfz��.�K�Er��qK_a���i!~�Żz�O=���A��w���� �Ł;�]�5>nv|�Sk���J��^5�FU	�����r�:�A$F0�V����8m�j-E:�?2#_,Tzة.�����|���kf89�0V)y�G�L��	&6]���u��|J��5���I�D-kO�֨6˕se�Q��3�3�%@�Qh�m.>?!K��ۘH,E�R&~�I�7�t(*�� ��`(�W�A#���v��R!RtY���X2�+�,<�H�F��݀�:�r� �t�B{'�\@	�=mR�F�>O�$f�I�rG[�ψ��BU��i�k�.��a�d�M�ý�X�p��<x~��Nd�9�9�}^m�Z��8S��L��
��q�,�A-�RyJ�0d�����N&)���ۻ&ɠ��)I�Q�����g]J�K�8h�b��=ǘ��g�.�D�>�j��s���Gŏ��U}	¸�����Y$r�5�צ��CH���:���{�x��P9^N��We������S�؂L܅�C4�������D��+����=inp���A�cn���?R�C2��\�H�o6l���8���2��)7�±S�"�gŷRҙ;�Dkh��u:���/Wb~�ntz����Q7��'����1��Ϣy�iW1�c-)�4��G/m��w�hC�oJ�g�{��I$�xqX��6������o�Xi��	bv�Jh:&�kb=b��L.�+2�*ʱ�0b�rp9��L`|C,I~�=YÚb�����!�I���/{et}N��v#�A鹼�1V��Ҟ;9�,�lA(�[����z�49���;.s&	G�αEZH�P#��|>��I�	J��G���& !�ǒ%։���S���?CB-K�Z�$Q'��f�p>(�ξ���Z �w7ðY�o �s��.*���|��Z��.�fEq�b �mqt��6�ZǧjO�A3w�1Ϙ�x�پ4o�M`��frf�'�{.t�*��9nG|8���k1<�{��P�]��}ˢq���:Ɓ�w�"@7�(��"ess���Z�3�u��C)U`^VIc	�rX����c`�k��� �#���[���(G�Q�M�o��$ʵ�^E{VcX4/.�gL�).���l�/��Ag�+��@=ߜz3
�?%l�Y�1���>�hl�r���_����S���a"6�7!9��xȼ��+2�v�4�pN�
 \�&�qC�v������d蟸��W��fD�C�h�Z.iN����8#�k[���h��
C�����-��oj�9 ����+�R��a����C�p��܈��Mm�j0k}���19�z)ba�[9Hj��Y�w���ܲ�)
�HY�+���^�tm[j-���)�-ʤ���c�@7�O4���qڲ���e�N#V��Ō��&�y�]���I��*}n�"Hbj�ʔu��z�Ch��e89ƂZj=�?�Β���/O�	%���/��0���$ݳ��g���'�5.�U��4�=Y���0�xk𹌰9x:�G�lD={꣒���*JZ�S]r]�g�M?EN}���3��k;�����O"x�t]�"4�
:q���" �o�s��޷�c:	��L��%�kW�������!}���r���atC����gz!�z�9�qD3t�NAY��`�9���n�vU��$�A&�q��{<��w�`��ŏ�N;����'�q��I�Y� �W��ޘ�zt1��:�	��!ˬ7�v1KD�H���zO�\�C��-��3G9.z�\��Od�|�n%o܍�T��n�� �Y�6!�m��c�^;�܉�NX�o~���t�Y �
>��J�]x\`��4�+����?}�E\�U�?G�\��3"��Y;3�)����R�@\� n[�Q���Z"�{��-�f8���W*�
v���sxԅ���	��$����0I1�R�z��e��1d��`h�Ё��#,���f��<͒���*#�䬻Kz���U�K�.��ʆ±��]	Jߠ}��Vd!Z- :>!#��.��+�
��d��>0T��)�R� <
I����G��*ӣ�֡�`�So�����h�@��kъ�+��C��wV�tf�M�:̬Q�Z��"���)�+pT���N,f;=�xJ�����1�@xl�%C?Q�(Z�#��LN����R��dP_��;�j��״�|H��o�`�efМ�
��������
2O_���:��ӫ�,p�IF��2G9���uɷ퍒�7a��H��#�(�Qa�h�e!��_r���]V���=��
9��_�n(�e�_o���F<�V'Q��p`~=6�S�DGEp��l�0�������L�U���oAs���N�>VW�S����ħ_u ���v��)C��[`��ㄴ�-��9�w��7�X/p�%.sdo�'hnK)v��4�]�xFe�?>p�w�;4��o��סc�̻����3�
~q�G�ᕀ '"�L����"YP8�ΚwNΠw���>K��/���E#�p��P;&���\z�4z�}�� ��zH��Д�)os�W^d�����ccpD}8�g��k;�u�dti�btxV����ܰ�a.����X�r*��%!�&�j�!�_Ł�;N����Y�_XtF	A�Ã���ZKW5P��am�'�i����&]Sz1���$=���vE�$S��je�;�8�����������][��^g~+�ft/2@�;�KrH=䇖��ɇ��Ҭf�.3������#N��L��A�ɭZ�dh.�+��>r�Y�J���E�I[Ha]�F��K�A�э9��E�[YG�O_��˶ON&�ڴpa�1I.�E�CX�5�LI#��M�M�R������O�!H:�b�B�|I��C�=gt�}'�g+�j.tzYM]�Q���2�6���̉W���|��c;ݬ��2 E�O�z���k��4�u�(�Γ���Q]eT������Z.m)~��������A��q�_@�F�+��C⽰5W���T���-N|�i��Iݖ������!`z �@�`�bb���V�}�u.Ĺ�c��0�&�j��72w{�0�j�lc4!�h]�ꪺ���_�����u�?�s:��N���w�r�ӏ�t��2֬��Ӥ��ؤgq������V?�9U�X|����^������f�7���XH7�����!��2�[�H�$n ��j���%U�� bc�Tu�huE~f3�������2@#�YM��=���������hv�����A=m�,#�Ge��0D�>��U�qn�3U��IXD@�#���FS�@���I��$��fbCP^r��+א�����K_E+��R�Z�:7���h����\�'S���X������
���o8
�)�@�3�!���I�x�G�pkIm(2���0�/�y��U�.*�NNֹ3�*�O��u�޲ ?_7���P�wf�G~�����"ް��p���c�Z�i:��~��$���ocXlxVHYEB    fa00    1500/�4��#O�\�Pք�+��r�PT϶]��6*�X�*����_�7vp�y�	�z�&},��_��F�;���-��LjisZ��o(`��
�b�Xی�+��Wog�+��;�֢��ٵ���E�@�C�0y����t�ܩC:��Jr�Ռ�_q��z�q�E��HGQ���7c��:�H� O\��n�ů]
f��D��|d���j�j�Y��!��1p��+��W(�NEj&T�B#Ηt��z�^4)�դd�1�DjbYF�������uSqÿP�ט?Da��0�k�e��L���kP��Ȑ��R�o�핌cb�N�{b㜫p���f�#:�9��FXձ�����~G���B �:���b�O�xMv�X�`���i����v���%j����=;m�qE�6��)'�a�F�.����	f3>ʜ�
l��Q�e]��f���7g��S#T�
���Q_��m3;�j��zu�e%�-v\��v�Y8Y��:������m�S3d>�4e @VS��g��q��4� x]/YnD� 7|.��r�&�� rN$ڂ	�}����D@*�iM�T�n��t&�C%΁!�"���a��L��9����ѭRV�3Y꾫5�E|&#s����=������A�PQ�?=E�bw� �臞$�q/���y&�5b�n33؇Hڟ��i��0@>Lj�׉�N�U�w�̶w��ͬt/�8r⼑� 7=�g��dC2�,�&����;�ZA�U�ؑ��a�,q>4�����]������{��
��n_�T���kF��d�K��V*�~A��$��3v�-��'��L�Fl����r��[0�̚�g�y^uwKO��n����@ɜ���!x���~�Y�Lv��fј��Njwj�ē�e�f��X=g;��G�|t���3J�O-k$/���x�uގ��nq����f�lw(��Qr��g.'g��﹮�|�9����*���%[�Ș�a�����1��5�u�O�M���M�+���hA��+!,F�[��+Bm�M�>Ӛ[����]Q��$/�(�7F�#�9�9Y�*|����;���Y9Mm{�=Ir����W>N5�Ow��ISԘ?t�1Znɂa��+]D�<���~0�sNݿ�8c�����s��2(�ʹ�x�B��/�ɹ��x;ል�k�&F�YM�d0���]D�����E���{˂��IUÑ�ʙJ���Ln���(U]��f]q&������t>��'��l�_��>ț|[E���١���pOP������;�)2*8�t4�=0�� %��TҢ��D¥��%�G���[�'uW�|��.���W��?�9�����q���i�k�V��󡙲G�D4
�{��ˏ�m�WL����!���N]��3q��O���
�m	yaK�U�����C���|cŶ���؉�������K<�[7�F(�V�~��b@[��<X������U�^-�iq��!�8��`*��L��W@�����?�B�7�w}�	E��� � ,���"$�Xy��en�1<��8��e;��jE�R��}�T^���KE�!a[��l��8��`�Bq���W�"�2k��{�&��Q2������$Ɠ�S�+�Q:m���h�>���T|�Ζ�ʞ	M���T��B�#�"ϧ�Yqm�B�n*�5�h{
%�t>��,0F��Y��_6f�Fף�}0�|5ý����.,��2���0F�&f���M����=\��Q3(�����hq�������2S��~ٴK]��Tʃ�^���[(�������W��H�2�����֩��1�$��J	e�����f��� 贪�����$�`������[���].qtAz�:�o�?r��&������D�E�V�Z�+D�87��ӹ�ɗ�4A(��dC��C �5���F [=A�V��`�$Aj�g |�;{m�l��L��-�M���OR$��ny,��K�\Z0}�_�A��Y3aV��;Hi�i&o�xm�G۴z?%O�9A�YM���N^�78"������`:�NQ}�A����)�m���J,z �Y~e}�TX�?�7�w$0}Ls_v�ܛ���h=���ͩ��%��6����;	=Td,?@|3x�����I�f��R'I�}����ͻ@t�T%��<�܌��9@e�u����4F�H�!	����l��h����~���s-��&���9'W*{�A;�d)b���[�I*ݎ��3yXq@�S��~��1A������7�w���ȳBE�>�/J��U%͏��CV��,����_�S��Î�i�I���BK;ǫU-�gK�"%���� ~a^s��n=F���mq����ԕ�h�y�V�kK�j��K��ٌ���}I��y�5�]kQ^עp�$�n�v��wlHC�����4�;? ��B�rk��YM�v��n�:��X�VXu�c:Њ"9�~�E�=�)���.]��
�����fǳ�A�g��#K� k|u�Ջ�@�!�+�3�R�[������E�)�l�1�筕*�0���"��S�����!jN��5_�{p���~,��xc�n���fY�"-���&_)ͪ���P�A-)��Q��gJߤ�Ey��Y�6UJ� ΩH57r"�:�WG��5-~�<Fe�h�1�bb��ƑF#1M�~9�����
"�� ���tr:�V�s�N ��6$�;����(��d}Eqt׏_:vag�e�oם��"K�����w�|ԛY_P��B�-�����r��A�8s+K���r�.�^nՑ��Τ��"�?�O��_`㭚Hj,����[c�A=,�'Җ*)����ϓ8`��O7����(!H��Utk3��6C}Ү/��ǭ�m)j�b�Wш�F���G>"7s����o��組O�����: ~uLx�ިz�WE#�����(�#���Z������Ij�x���t��,�)��x5��?�EJ �bmZ�k�ڂ�!'��3��R�A����u�C=�m2*(�5X5�v^�R��/�WP��LНm��J^>��=���OE��G����}���MEɖf�M_$ �UTc!;�K_+Y/�>mK�v ��Bng��]3
K���'�|��4�4F�r��5�ܥ��g��Y����_�p$��k��f(�Kn�� �fܦ�]�$���4�o���ϗS���J�-W��ڽ�V�/'v��f.}p�ĩ��s��@���}��^�ft�#Y���U!�¬W���5J.�ܶ�v�j+�t�'ޠ���|z
h<XT�#���.����Y�����={pLr��	�̽������٫��G�_��-�r�����Eez��Ci�}/j�XD��1ЌNk%�p=U�ҡ�9��%��{ �pI��E\Z$�� ����8���<"s��UN�[e�(�O�ނy���3k+2�[�=w=���؋.����8:��뛾����u�	�Pq^r\����Eݦ��f�p�  ��"��{�4� `s��Ȇ��Ad2�|r�۩~ ��D������t%(��%�֗��߉$ɸ
X��pOD���(T���	 7��ˌC��Ym9��N�f��ɪp7�܅�/���?�!x	1��p��f��y�w?]�.��虑�|�ۧ�O\t����ם�JG޵�ع���Δ�o)�Q'�s��M�|Y�ŗ�s˽/!�/�G�o%��|��^}|�O�u�p&5)��ͦ�&HM��T�5���r���Ǔ�I�*�u��9&�J�&��w��I)ŽK����e�է��`�*!7��ˠ5������d�C}���y�#4�Z�ˢ(�4����8KP��^phhV������K[ٌ/ڜ⧜Q}y�N�$N��F0i]i0����z��!�9��K�Wt��NX��]��,�����/�i�����p�'Ա��?�/������a�y"_&u�K� �P���n�	Ƭ�HsыA�n�J�s�9�eT������lyH2\��ƌ�N��+�����T��q[ę���{�Ɋ����k��2�����-F�۬B:m�W����N��ՕiFlmrL��Z��AC���yFܮ�L�(�*bS$)�k�;������,�6%��W�֗�Hx�i�Q��8�������n�����L�qʊ�x��~�O�v	ehߊ���2���'�� �����v�$�^AK���f];W9��L1�����Ѣ�d�	�]ŕ�GZC߯�CbQ�M���FI�Koڤ�z˪QۀZ�6�8"����6��	���ɛP4h����Y��=u�����<]��w�P�����D���r�DE����Kr��ɉ^��r1�O&�p�MoP����0���_4�&|?2 n��b�r�%W��7Č?I1#mӁܓ���+S��0��J�����D���D�~�m�K"X��c�w��Oث��X��z�W�
{�����3x`���ؕ�W�Rꗄv��.%�f\όQ:Ӕ�[2a�π���g?=e*,]G��R�˄(�~�2�]�f�R�^z�d��7�x�8�>8�}�2�6 �Y����[��~j&�֔��@H��/
�����)e#E��e+��3md�\��aü^w��J�%�d ���o���ؕ�L��y��U���%����w85�jpKS�  � ]D�7µ-V+0j��i-���`���G��ϗ@�#����r����7�!`�=�?H�d�G��\�&��|��6�9a(��
<:�I����+7��gq�+�+�T{M�xD�1bi�xa��RQ�+�����=�x�^�y����ؑO]J{��ji�x9u }&(k������,����'fW-�`�<���k�Mm`��_��z��E�$ՃpR�[-�����<��i��.�!�jŉ1Z�,���2r�9�\�w�+���#����Q;�f��L���iLi�m -D���S;{��M��g�gR?Q�a��4�61��)E
�gp�؍L���ņ���@����`e�ތ~���GS) ��@��!�{j2���H�b���;��g�\���ǹG��Y[g�d��#�-z�9`42�����@t�������amUz�dW�.O��&s��"�52�(����e�`~t�Jw"j�7z�R����g�Y@���w���U���Yx�<�
.�\Y$FID�I���!��u��;�}.�mA���S�Y*���F"����͹y!.ɾYO�K���[f��R�2 �{��[�3 U����;�/()5���M\Y۟�m67�����jw�[XlxVHYEB    fa00    16c0=_T�MMok���`Ӵ�5K�5��(XDC�m3Q%m��i���I0#���϶���0���܊�x�Q{m��FR�uْ�%/���w� ,OԒG�>���r�y9�_��`�����	y.��JH�cخ�*�
�'ҷ�X���%q��B4}��������2���.���z�ܣi��0c�e��W\�2Sf]������=�Wn��Pe��Ì�W�Bd��k\�3��K� �x4���y
R��)� K��ڈ������}�10���T����7����{��n-BZ���9�7�jI U�:kK�q�>���T%9fi\��jF㷕��Z�O���:2u���/��B������U�0�V��]���sC�U�x���I��,��8I|�d;�ʐ,�[�:��h��gZ�ۘl�%z��\P���PԿ�$���m����>jB����G��\���w tr��(��.T�R/T�`�n	|���o������V�wzև�K���x��t�w�E���?�Ț#���}� cc���8��(l�����64������IJ�p	]��}cu��Ug�|#ID��$K���r�bB��G��h���T,���&����9���?���2��!�+�~?�N�oӬ��ྥ�L��Nۻ���Z6���F���S8h�s�Vd�p��J��WJ��j��g�<�:��I�$��F��X�qT>Wɇ�V��m���@\��Q�h� Хvp&��}��g�B����8+�BX���`F���HM�ce���t|��.�"R�,���}�^[@�5Z�M.�� �EJ�	jg�����;l�9Eg�8v;��4%�sdwi��0�}~��`����Q�*W���NL����o0]�"T�w��@�y�v��q�d%L�&qF,W���U��s��Xl/�폰|+�u]�F�V���j���=NK{���J�~�zW�A������ck���vm�ߍlSo_��tH�h�����-cpb�?�3*ۆ�C=ѫ��W���J��{�3%��Z
�A��t��w:��J���w����K�n�@��PF/Y��o�*�1@���n]�z�Ot�'����FE� �AMSD+:�x�*�$Ѱ�>!�Ѩa����F���=z��o�:����6Y+م�B�,L�T�K7�y~�͎��S��W�z��֣
��q���?i.v�s��؏I]x�� �rÂ���b���C�O6s�-N�����b�Ѻ����%ƞ���d~����dCL�]/�Q��J���VQ<΀�MIQ�K�2&��ڧ�$���1N�N�0kF���b3삭����h�	0�^�V%��o���mE���-te�O"��D>a�ͦ�>��2	n�x�̈��X+(G�#)��Y.6��q��ˈ� mа�A�<�:KU9��".�� �-�P��Vc��ؙ�K�X������O
c��M�s���U�;*��Q��_�NE�T�z���c�@��Z$\5(9��៯n�.#�o��״�������ڕp�XZ+���o	5���){z�:��[Z���r|�]�&��z �E�侦��usׯ��eT��t+�U�*~ݫ���8�y�ЯQ9� ����V�N��_�	N�*� �e��a�_+s�,��;VB���p�	���IVZY5'v����8��v&���<�q~"�Pr&�xQf��� �-n������S�ӒL.V��zz���l���c#{�$���Ϗ|�TNd�-��g=�S�.�ȍ0�!�
:��&����~�}n=l��8n�E[;��
}���f}�S�V��B�,�Cߢ]t�e��>h��J�
�F����c��9�
ˌ��>'?�,^�eߖT�ݹKALX-n4��"�b�H,,^��nxh��xk1�A�,��Io���'�-2�[}#{�3Q�@i����O�|=�x��[�\��#��ܶ��r������;ks{(P��%HҀ��Y�`'���]�nl.��DLR��wVLA��'{��v��<����*�ʬ@�]�nfL/Xdͮ��5�Nͦ�V����'=/��kiWBѓ�J�:�bKu�^l�q��k%��{_ڱ�+�C�4�6�Xi������mѱ�sH�J��'��p3�MdkYUN������)l�͍�,[�����6�Zɾw}N�Un�qPF�-C��Ԉe
�'�Ь�<9N�h��3��nߟ���x������Am8S�/Wx_����_һ	�)����Y����0*-us�	+*�Px�~���A ��D��V��`�
��Y'e7&�W�A��ו.9A�����CkI���N˸?C�%�e�h� �C�L&�eJ 8���P,ě��4�B/}�\S�r]�/G���\gv�ص?1�� נ�WG��n�U� �(��5}��{���@+�eE�Y*6/�� ��yT�i�T3Nb�$�P|`�#��׈l�a�b�B2@�L�pŭ��	��{����;y���3Z�?����Ł�M�=�3�āUmCbp��A�پ�ũBC`�" ���#)��O]�o�öX/Çش�����
-8�-n;�B��@8�U�[��P�������'�13O�LE�4�f�߱ij�!����ov���3�(�za_RL����J+�}B�W�!���	,{W>�c�`\&k�ߧy+�tB���/J4���X�Z�ugua=�s�XFQ%j�4��io${��m�i�;/U�M�����������4x����ϭ�I_m�|��3�ԫ�s����Y�L"7�Q�X�WYIJ�nA� ���}�o��	[�Y������������	�6Q�,�J��R�iS�o��Oڲ3��ˢZ�aV�0����\���ػ����1��Vb
_���\���LH6Î"���<'P!�cF�=r����'���F��Em6�$ej�m?��� �ԧ��T�K��nU�m[�S�f%ѵG��F-���[����~v��b�k���]n��)U�Bl`Ճ���j��P����b;��A*��HP�t��r�U��i�9�:�/U�>� ��R�#�ŭtM�~u2����`���~�'��&ŎX��3c�ܕ)~0ueikϤcJ!r@n;��12���M���w�/c�K�wxV�շ��ㅖ��i�_F-�LZ�`�=���8�
�*O�QSwc�d(@�#`�=��]
&�r����srR{Tq���uD�"/ɳg*���2�p)8ʄ��V%��:��b�/Y�`609���~��z�"�Q,���B�~(���d�r���<s�E�Y����b;�y�%����^g�5+a^��U*��S襽~@=Խ�_8���a�<�R=���<����j-�"py����?c)7Sv�'�ct�R,Uh�o���g����*ϒ��X)�4���=��l�h\O��M�/�\e��]�(��T��ʮ��z� ﳊc�z;�r'��/��AhG�Na�4Hl���I���?�����N�G,���G}U��@���e�
]"����P~���*?�Z�dj*�"4��"~�������8����<C�1WUD������ʄ.��sw���e���.��,!�gp`�#M��12
�
�vJ����@�T?�j���!\��lѨ���b�ⱅ��õ�\�M��͡No�y2��v�o��NO
?vi�BѽZ\���f�i��� Ѭ��Ut���%
o?,Mg���W�ڂL}�uq�����vzJ�\��p�z0W6.�oٽݞ����HWt�QK���I@i.lv��J��D{������q	�e;��c�pX7���zu������'�l��v���Q�ѿ4�,�A0xω'|q���jڗ�w�XV&k���B��qYfZ�~xo.%�.|�w[���z�O�k��i��g�(~��`�P;(*�Z^k�X��"����ug(=YB�:�$� �0�3P�*d3ށ���fD�������u�T/��>���ky��Z�%��}��d˙Џ #kC���V�*+�L��7ԝ�7��R5lY��6-����㭮�����Vay8җ��T�eQ����Y;N<�ϻI�WˑZ�/�y\O���.���'EV�}�F��g������!))�#t�AT��ƻtֶb��� g�"�c�?ln�_Rtf���e�z����I��
��r��]��mnT��S�U6|$��a
=���EKrM�+:�����b
s�a��C�[����ܠ(��~1�Tlre[|��Ƶi3�M��쑒N�U���Hs���-�SF��?	�`� l�ڻ#+Y� oq��_N�KꠇH�����A�E:h%-͊��/-Z������X�c�m�`Z��9&������9 ��+<��H����8[(1f�O��:��	AT���K\.��\�܂��T��ؒQ5
�J���f�M*N�{���=��k����鷪}��R���,Nߘ���W�F�o�lB�7�X��kF�J��K���ثV�����R����rŹ��zC��i��卄��^呹8s��c�i;��un����i��[P�.K�@�2�O�]����'-�{XS����?�ʞ��� �e��0��!s E)��Q�o��kj�^�/a��h�����J�f�qD�A|>J���(깳F���>����{�:SM��m�m�h�t�ЀV$�Z�y��/:���[��HBzW~>?W�nź�)ꅙ/iηp�T�3��#AMz0�|K�1t�Dևv���C詝��� !&˟����˅�p�;�2��T��U��O0�Fm��!ͺ?'F9����2((=;@� Mq6�zҩ�MG3i����'�rDOI%!dL�7���pC|^��8�Dc�ɓ\r���޷�W|x@���ߏ*��b�L���=�7�ô�$�{k��ٻ7��J�3��&M�f8q��:�S��Ld��������IE�CR
����{:�#�CἙZ��cv"�0@�9�ȱ�b�^*��}`��A�3�<�� -�!p/�� 7�4��Q�dL���j��v*r'�A�_Hn��d̀� ݱ��o�sf�{GVr;R���U}�����T����ޮŅ�gD��^=��Y�̺h�d.H���.�$���	eq���_���,0n��"�
n#��?U���H����ETYiY�{[��X��L��	�t%�s��07fxk��āI�kY�2�A��[�����ؓ*�ކ���w��$XF
�b�����j.�f�A�D�Щ��@)+��ӻQl�l�4��t���E��J���1%Y�P���͹{ɮ�l����V,��o�}u�f�?A�s�t��Hc���G6�[�.�A�7Q�h��;%���n�+��nK�e�ϒth��!n���LJ�o��I;"ʮ!����o�n�,�S��o�}ܟ^b�X�#&��`��8E���Ȣ'Bf,d�0�ɫ�~(9�"+���(\�!_C�d�����ڔ�G#ty�������uj��T&��)�}fR�����?��k
�љ�sz{�}3c���9�x¤M-1A���dKN���H��Y01�K����&r�`����w0����_'Ѹﳉc��0C��D
�/�&�UW	JA�&<��F++���0S� �E��UoVKXin��)�9���B�'��^���	�G6�}S�ʣd�� <-څFw�L�|E�6?�XlxVHYEB    fa00    1740o^�rRa��A(������I940sR�)Z������������A" <��z:�`�	L�HYH[j?'������o��:�7]� =��!�|�����A=�yإ�Z7�U�%�.�J\�/��;z֌��H'��+�g�"V�Gr�\��z�W�?��@��tA߾�����Y�����:��Z$�H�h���4ǔ!�Z~���'sd�����z��郒S�;3hk���.�NB��O�a��e!����/-��=iY����'��<�/O���:5*K���7�Ֆ��f��S2Z�����:<��r�>qS"�M��S���o
.��*�2>HAK��v_RY�R4G��2��ʁ@[�x$@7�t��N�Gy�g�M�����6UE�^ ����D ���%s��e)���_�-�f��pƹ'�w����P�l��GL���~-W�W.��cmhP�,�
&F��	�G9E�șz��b���/��2{�9���&�G��'Y&4�,�'d�i��@�}�<���B���$ ܑ��;�~������_nVv_��_����C#��Ғ��&������K	��)X�.��;x���(�F�E%�*c_'A��q΀VĨ#6sH4O+��!���~
��#�ϲ҅$��Q4'�Ȗ�����\�W�x�C��N7	N�RԢ7_�R(Њ|H"/�LJ��˗��Rb 9�pK���L\RC��H�E��Xa�}�[���Of:�<~�BYO��mbEe�-��j�%	{�"�@ps7�uT���n���\}�~��F��@�1��93��xT��\ͽeZ�I�q�@*!*�:��ό?�+E�������D *�a����l�Ջ��cE;Y?��c�e7�V�#fE�_�!��Y�8ߣn���(�r=��[�I.Gh��
�-����nb�ffn�@��/���/��t�靦�-�+YQE�	�)L��P;X�6 �����iY��I�������v��,{�$ƹP`��z��~<����?vŽ��os�凃@���И�RjǙ2��{@l���Q�����iy�}s����=����'�����a�^�����y�<DdL�1����m����ᤌ��C�\3#D׌FEN���w#�SeK5�����^�Gl$�� W��,Ȏ���H���.��`��	OjV�W�
�i+�=wQ����� $O���C�Yx�,+y<3�8Bh�����ZG$uG��N:髷RCi��;pF��(�C<2���'�� �$#_X����� �<[�p�e���������q��R�W��X��dyD���Yy�U`��x��w�����u6��z@�*�eܵ�G�O�+���i�1H�:��FaN��3`IbЫ��JV��K+yޜ���S�t�V�����
�z,���B�{5���i��Oݻ*΋!��=!��մ�8�!��LdpV"�
�nvfN9�<�#7��m�N.�6F'!$|}�?o0{X�Or+#rE=�:����UI$鲁}��eZdѲ�0�-'5k�GiQV�,��o�%�F� ������ԃ��P����t��4�?>R)DJ'� +nRav�qV%�;� ���z�v��`���@9���b�p���FVkN����i��O��П'%P/�L�4���b*Lºk�L
��3�����ń0뿕�_�_�+c�x�¿,�Wa}E�Q��}Q7 �';���\f�̕Ev>���cq���Ξ�Y����dS���	?�Og��y�7Zy�˭�Q�Vpn_��j�*/j:�-G��a�h��zQ~}�-�d���(UY��O&�H�p �z��l˕���Y���,�7�d��;n��� l�I<@L���7���R�8��Xj&Y��1RvޑM��8��]�$p'f�b�U��k�EY���v����F��F ��؞�إ�l��r����܀�c �x]��R�#��ʽ1x��~��D���uE���^8��t��mN�թY�0�S� _x`G [r�q��V�WUB��gȚ�Pm�����D�cɥ�n�e�D�I��b̬ B�O�
HI����)L����%	�T��'�cw�1�����\�c���`Kj�<��e#��ss���?5S���:�`n�� K��E�)9/�f�e�j6"��ZZ������C�"�R����մ�CP��|_i�"���q4Hs�[ʂMu��!���S�H���Wԧ�5�2�b�w�ѳ*�4 <��ߤ����E�-#���jk��ʁ��3�F��\�@oj���9�f8�����EiwX�sJ5��"��K��د~AE.y.�x��qR=�� �`1@GQ�:y��Mp�����m%�U ��C�g%��AC/m�k%h~~f��ϱ7D���2�LC,�m���*&u���������DO���[��`���2���c�v��g!S�wu$���T��k�l�lٿ�S���lرVd	�� ���D� =܌m��
x�QU�,lk%~��DR��[�!�0�籋d{�@\��~�.�h�5<��L+&��T*���;�m��Ek�h���nqT�BL�t��9��b�r�kw����<Y_tUl�w��9fT��ӟ����$�R.���˃桕}��mv��Y���Hq�9�Q�C7~�얿�T.^�E�?��<J�1Q:��j �ڽ VRmi<���J!���.ŅWgÆ��V(��f1��<{�"�7P�8�lWþ�K�O�)�'��b:�#��1���mo�nF�{�'���sa�=���JfD��!�>�)׺�w1�O�>Pn[�3��4��7KM�����%[7�O�Lv~�4!:Ah��(�7e4a�����*�>����5M�Z�V��b^��K}甂��n+��y�^���F��P8��ħQX��Y�<J����x�|}"�@���8��B���^���0c�ouۼ�K.�T��R�L���j���޼�gp\���;�2C��պ6R��F�Y}{i���V�u�ͼ�����sĲ�5���2��4Ռ��,t��Ȧ��+!Z[W9Į)d���W{}e����� )u�A��"�}ѨM�NHh�3��z*�!U+�T�
䃠�9��<��@�
���y�z?sW�����W�I���������cg��
�D�@K�sy|w�	�$r裢^��f& ����̷�2*��)9�3c�q��x��p�X� �t�@�He�"a�Z�Q��`�E�vVĝ���s��m�ZE��yS�Z͢��8-��"e�F�\}j�
�5���5m�BGB%�`'���;ꈍ �����	��`%�f�D���7��H(�]�W>�I�>ͻֵ���q��W��ʐ�2�B"
2b߫�p8��jM|.���Ҝ��	�����}�2.ߏ|}Hm|	�8e�����gr_�)�r��ф��Ys6dU�T�6f9�>�ԐsN=}�����_K��>v���!�i�=`�+��6�2)h��ǌ�C����wv���F��aM�Iq^�$"q\�H��x�T�Gn>�e|dit�V�*L����p�gG���E,N�t��.�����O���H��R#Z��<R@y2���pgsU��.�e�_%�������&��t���F,{�_m���\_�ʇS���1��̡��{��Y|��i�kٍ��@l�?1����wD��C�����N����Uo����ULe��'�I�H	�T�K��l����&��j���x�V�V���\{�x: {81?�&L��e'��P+�{nlJu�f5	�eYe�6I*��,E�ח���]Z~y{,�ڐo�+i�v�l�R:�K9f�����חUyRp�uLڮɷP3�u
~�����)I�F���-�3�b"�b'1��X��� ����Ⲏ�gN�_O9C��_V>�NݝY�V�SH���OdB�aI�*!��`5Eo
K&\�����
���`ޙ�or��h´�Z�]7�>Dj��%`�.5Ϭ��I¥����>�>9;�	�r-���
��}�"��}9L�7D͑�ڏ	�N�Z5����V�O6�=ZO�?��˃���	yLmV�v_��S���Q�&��_��Zaꝲ�����lXēx���`���Y���`�w/!��v�
��1�u�~��.��� 6z����#�L�e�×�)���t���l=�퉕�Z��B�La�k�d>F��4z�%�z��lx$�#��g�A3S��r��Jb�"���n��2�a�>c$0ƾ�y8�"d�7&Ll��w.�K8HrZ�$����V�9�B#����b�[�`,=U2��|^�.��-�a��Y�Ge�;�aQ�^sf��킆�{1��հь���
�O>��C��d�R?�P���p��GR�)N��պ+�0�� �xp�����e
m������nM�D�3�D�o!K�,�h4�ሂ܄�;"�v�#\ϸ���9�����D[�Q2��M�]�c�m@lJi����\�g&����^�t���'#BB�P����5�1`��EE̖�ztb���rM��'���g0%�`�ג=����>��Z�;�����>�����C&���t���C��B�}�d�ۿ��?��,>���F&$7�AY�]S3��z�+V��T`\G��p?��s�
�I"�_�w�J�
��'�G~���C�"a������!m2ۨ7�O��&b����� NTW��j�Qrx����Vi7t0�};4���"d�=`	{$;d4|8���E� �\�+��:�V-��b���X�q�f�t��:b˂(����<�����8���A��N���)u8D�$Т��ԳRI�2�5Gb�Q�)U;�����6F�M"H�<J]�<X\K��|\d\`�y
0�= }�+l�=I,׵��/iB!��ڊW^�u�}�a�&xƦP��:�ۏ��$%�Pڸ�\Tik��1+O7�`��rى���t�o4T���lOp��UL��Bv	Z3�)�c�gr��r�i7�%K$a�V�A�+�r:³~��o�^z!�u�+��.��������w:N�?��v���7r"G���]j~l)�ں�}����-�{�Ţ�ԿSKg��6�����i'ܻb�
_��~��&�*:�M��C^�/rZN�GsiV�g�_&~vG^�#�v�p1W}�(�?��/�<����M�P�ё���S)3�o��׀�ke�0Z��\b�'���5ڠ�{�}���L�o��qnPZ�#�~nU\���|���e������>/@+����h�Ԫ�j��G����n�Ј Ȯ gc�Y�t;:�}l�n��c^l�۱R�b�wK!d��D:DK�l�`=/\3o5���7f ��m���dq�h�	����[��i��6}w� _FD���w
�$����!�1��^���:�{����I��������oj]�����k�8�1�Z��x�[+D�B|��d��X�8[�6�P�I7��/��(&���H43������Y�c���?�1x/�O���^qi#�^<&]�JKf�;L;v������}��D*�`���0ʒ�+r��}��),����W3����� 3�\���"g����u:��i�AX{��1@�I���
<r�I <t:>S@؛j����]���c_̬������'o6Hu9T�D�G��d55M��L�6��n(K�Z��Z\�ẋ�N���E��p7?���l/P1�n0�+O%�(��er̻\�w-�ːȆ�Z�:��=�v�Z7z0��A�C�tPdNr;sI��e5�s�⼛���i���P���:�>�m&�c� �#��Nп�!j��O9ʃC�M#G&�W��&�cJ�]GX��o�?�u 3bM�~�J4<SAܸ�lP�mn�����D:��'�*8��Zn��	XlxVHYEB    bf14     c60�!ey@�]ڻn��u?������4y�)���pYk�b!Y�=�˟��6;�S��cx�3!�Pw�L����>e��M�?�)�
����	�1v,�hXބj�6�o�K-J�}W�A���.Ϲ��VѾ��-Z 0��U@��k0�t�k�/�3(��@�.4%K`��.����O*��{{3�~˝�4۷������V+��S�a3-�;E�����	г(����%�{�2��"�;S��{����K�Q����{�^_`�c�v�l���Z�}���WK
@j�}ة��ë�{�(}Ҿ�k���d�h6�Z�l��h��on�ӏS{���68�&o�{��
���5�J�2qNU}45�8uVV�h���v���(X.���e�7L�45����<�疉���1n�4�lsQ
1����_�E�h�𛏧�\4s��S�s�
�nq�M=	�8&B �k�B�;$6�_jv ��K:p�P�c�]n1��R�Xm~�u$6$Z-��H�H݇bō�O���>��N�סgj�|p6����d�0xd������x͆-�}�sk&8~D�4�MMA+B�G�wT�,O���ΌtkZF6��0֊���}����e�������"�I� �:/r�$�F�C���f&���H���\ԣ�$��r5�SAv�����'
�B��S��]��vZ��ʲ���Da2�%3u1��M�L��q�>�0�m�!�-$�x��ʍ~H��d�h����^�例y�,0�7�
ocE�D�� �/��鋒\|*�D�{y�ˏ�5��E���g��|�Ʌ�ah��I�zէU��c��Qs�[��q����)^�J��Q���	��LO���	x�w�"�k2��C�!P�`O���{��%���I5g_�f/��WQ-�h 6���S�O��a��r�tP�S��UY/7�p��f�5`������<"<�֘ng�R27xs��)V'�7��&E�+f�|2 �j�_�e��Р�*�k!$�:e�3]�`F�L�h�#�/1u�B�d#�`�XOu���ĝi�q6�5�%����%Y��E�VoHG;&��Py#oFz#���g3�Kb�%����l3� �����T�ƕLBZ�W�R�r����<4�lȃQ�6���/�������^q�]Lҭ��sd�a~��!e9��{�(��F�M�l�����C���k���-�NI!<��y��@8���������Y߯��v�|Z��K�^��������U�X�k�3�Z)9�$�h�*��`��Dmr^l�ge#[Pu�e�^.�ɿ=?dha���D���"���8��.\?T��*�Y�NKr@�C��]�'�|U�O
/��a]ߪQ��,�a.
A��������r�l	݊��6����ݪ�c�]��]���H�ߴ�N��䞸��٧�7�L������_ï�����ZL�؋���)����c��t-�ksy���H%��u�th0��eη�P���M$��ǵ�;��{���n����{#}�>�Abxs�&2�3�C��c��RË����KK�Mf�
���*��5c�P���p������nO��OAѼjT'w�����±մۑ,؎���;��q��,����v��P�VR��r�z j�/�������ı���̀��o]l���ؠ<򑉋�.sq����w��S�S杽ݷ5��_��HA��T�骑��p�V��dyp+��;)���Oe�m}��
w�;�Lr�Q�^�U�5�]S���샫�z�|l���x2�\���d�v*��َQ?-��r���S��_I,���%��ܚ)$R�NE�۩��R~ͣ��
b�c0�X��G�<�䷍��q�3��w^ ��U�C�S��q%%v������6E8r�����Bي<GS�L���M��jQ�H��&�`F�Y(b�Q����?"Q��,��PےƣmmǊj_1W�, ��u����E�(^��Ya��=�Hp~KH���bJ���۪2D8��	^c��[J�����_p�ZG�Z*Ǒ1���e���Z��mЇ�i�������%'R�h�2ۓf2�c3����>�{eO�_{@�_�Jl3�+ឡ�������)��[�]�ur1�C�5
o<"S��yY���M홳����E�<��>���[~��"�e˝�=�AfV�Cyq��\�6�|~��c���T��إæht��#ͣ.	�����0���1��;ȍ��ݦ��<�M��ߜ�0���Q�ad��,�~��<�[��B+�2��������g��	[t^\��*	+`6D&S:}�Gw��#3��F:l ך�G2
�%��ڷt�am�������f�
,��swѼd�`�d�,V׾��Ӹ�;�k�.J�%LRMa@?6j�zU��WS/mLj���g���^�$8��F���p�?[�b��NKQh��hgƦ�ɉ��lޘ/���k�)<r�`.sv�W����H։{�����մ���z�kUx%�	��+N����LKh-�b?r�"%����[����s�yn����[D�.������K)ŉ��[��̀CVT �Z�m�[�ʁ[*}8�Ml����qG\x�P��*G0��i>�D�#�~���(Fy���Ѥ���P��հj�iQ�V0����R��3��L˥@�cJs��㎐O��������-�g���֦2#�������C�G���n<|����ÅnDki�i�֯��֭*�>�"��4+�#�Cr�wH�F�6�?�E20-�11�Jŏ���#Ҁ'*�5�$lv��O��)��rO���wa��h�U$;0y!������׭=(b_2Ș�q�e��0�T,�;�QG�\�7W�ˉ������Ùm��l�V���;C$;��t�Z��7d�t��@�ї)� ���2u�����YPŸ����T�;�EDԻ���*����(?�qGOB�I���Ft'�Pg��}%xخy��~�#�����s/ �~�ڻ4���o����̖�Z��"@m��~���`�����vn�J9����z\��as�c4���J�����9�rS�_�0��O@�{�_V�����[j�!�f�>G;����U{"l�Y��