XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����AD�h)k�K$��jXxu���9�b`��Hg���(����hX %N�O�U;,���n��:�)s3��^g� �Z���m̟�p�б%�8� +�x�O7�����*䝝 +f� �x�4����QPo%���E���2[�#5֒�0,!�[m*��8=����G��Q�
�}��2ܾ���c9zd��bDO�*{��6�.f��^2n��4m7�R5E��9�ܕ��lв/$q�D��CD)��ܟ��8��v�hԪ|�R;j�aXlR�7P.��ҎM����~�W ����.i|��kNĄ��˶�-��u+R���P����46z+ֿ�D`��b|���S!��+R��_��սXp��ݙU�W���P�M
/)�0���9�5�l4/�,%�E��J�9�L��k3�bC�.Wn�m��A�Nhg\�8D�5O\�UV.K�:{�xaRJm�Ո���́�Q��q���N�@z X��!.��V(DO�%ӫ,�k �-���x��l�)m$y߶��S#a-�P(	��,9���x�n	Hk$V*k���;n��?5=�qd�7k,�:q��Jk����(3(���=u�c7g\�.�^����_�,Y<|�'���B�&w|�]13F͟dp
�x�"^��g(V�k[��:�f�t�����7_\�>����p֢�Hvw��4T8�b��eT�,�ȅ���P���~hd�(0����meA����b��8���v5T �?��"'z�Eu`˖�>XlxVHYEB    fa00    1ca0ź�*��^��z��#�9�p2�w�ޖT9����Np�ej�7�"���Ü�bBR���7^H'�t��Oja�������3�� T��տ�\%�v׻��
��"�Q�p��P����/������,���X-��e�S��ɳ�
(Z��)�f�@&�B����|��vĔ��@����f%���;�7���_E��:�OLҚ�?�jj�:Ԧ���*�F����Q�tsh�سsB�������:yZW6� A"Y%<�8v�S��
�!k�D�~>��W<�%�7����ru|i\nhJ�z۪6M��C�G�GЁu%��R�iu�g[� qGg4f���	 u�&ɸ���}�-�<��-/���A@��U0�p�w�ӊ4,�<��xI�Ir���Ēg_{O8S9:�q7?%&9�Z��IQ�o�,Be���Y��-Y@���[7�t)�5�{6��n\4za�w�K)I�0=G���Z�e�$P��dK�*��ں�sw��P�Dd5p{�T���#l��&�t}���L�J��Xq<�8�^���.B`�Q|�1�ð�q���$lI�D$������â ,>�<-љ�A�Z�&�:������xD;4�q"�,L�����k�iB���>c�O��1�����T�Q��Z��L��B�����ˤ��ʃ�`p	6�U�<l�\	Sɰ�P���kp��T��>�;�$���θ�f{�y�qk{����m0:��(�7�bm�Q�XY�1����[b�����@R�l�
s?����8�p
������� W82���U�]P�~1z<�Q��t[�"�q�N��N�&��YhX!?�z~�?���}^�9#�����DI��'��!�O4X�_��c���bQ��_��6�a�@��� ]��d)b���i=��q�{x{���謭dlT/.0�3��Ӛ���T=en\�X9_�/���2���	��\DHU �4!_[g%X9��u��\�6�}�S���@��ln�O�S|J�հ��C�>b��|r����g��uЫ)�3��!	�T���XOq���єQ�+&��G��k!�ϑ�&Ok�K0�E,��R�Ng�Y[D��WS9�V�z$L^�4��{ehv��	MvK�D�g�}lw�u����{d��2�vB���<ο�;Efʬ��	����@>>	`S������e�3��p�B�0����ʪ��m��O��"��� 
àK�(v���'���c�+�M7h�!lʆ`��1v��C�8��e�c�m�ӕ�wLҊ��/&!'���:��m��v�n������N��yg�͜�%�j�Cn�_pF+���w��Xp?��^���-��Q�;�k��G�{�M���O�����$���Z��)6DZ84-e�ݚ/[�q)�؋���p�<܆�|�Ć��	��s��9*��i���)������G$�O�5�O���]A��20�����2�PRیZ���w�Ⱥ�+���+t�q��;a�m�	��N�"/�j��E~�����lDSQ�}����c�L7K�v�t���e2@L]�B�,�����߫lZ�[��^4KC�2�с�#���E����K	�H�8�}&P4�-'�k��7� 1����r���*�(?4u6��n�Tl�e�-��w�'�nvx����p����x5^�9u�	yT4s��4��R^��qi�j����>��,�ۚ���|�����Ϸ�.ohvڻ*UT��H�g���d'���E.���h��Z��#+[
���y^�{K���&"�����(�(�c���)Ĉr��HYB�8U��E�%L6�֒��"�J���U�$��c��+]��L�|��d������I��s�#������r�ty�m9�g�l�p�g��s�9��]����FU��%D=�/{jJ����df+��5EElD�٥��������2�$����?��x�����#ne7�19��K&&��� ��#E�1���X.�5�I��aS �;H�����������X鈂Yө�)-$���+�����1��	�[��4u��ׄG)�[x6�+�y�x;l��0w���=n��Rw�j0<�r<��֎t��-5�E�������̴Flo�ٔ�g�Gf]�[�7�yq�c���
�cn��$��i�(�%�qfJ�|��5Y �}�g������0�I�0-���8|8���!�-�UFu�H�����C��G8<[����	���5&2�Q�G��!�i꽓�1�b�SD�y��%2�>�) ���e�ώ��{�%8��4RY(c��Q*I�YY�P1�`�X�p����s�%0 &��?�g�6R�!�^,F!6ǔ��Sww��� -�Z24�7����l�l�'H��˝�q�n�G��r�p�<�sd_ok@��H�����M��Q�¢���e���sd����
��ۭ~��>�L���jl�2kU�9m�W���|�[��@�(�������K����L�C9��J��g�M���0���z���N���[d^)ʼc�A���T�u�jz�r&_�������x�ZUӸ�u'�M?�{ �x=eDAU@�9T����䬾D��CA�4 Z��+�!R� �o�����������%w=i������Zc������y�� jz�'������d/3�saz��SU"�۶<���ܒ	�5˗�s��_3`qc�/>bly��|l�<��mf�쉓�Ŷ��WkA��2YsXt��	�U�;#I� �-}:�;�ǭ��֌a"۹��P����©�b��뎫�>`ܸ�[s�I!�7wj.��M �jt�gYlCiVUi�2'c�cE�(,{���6�k<�I�G�g]��9M�ܗ1=�H����3]V�"%t�x2t�H�w7�pɺ��N�(B)�op����6��A<W���J>A��S ��N�L�2_���f}5|���V�Fmc�g��	���B>]��m+���&�qͩɊ��_�w]YM]��B���X��@Xo(��86�S��Ѻ��L�]�������v��)�W��f�f,���ZVQ�Lp��D���T�34�\���@�quxet�P7�	�&�h1l�4-�yg0��d�Q��o�r���]�����muJ~�[S�~
�z<�$z�����oH��>��"VU�f(������q ^���AM�}�����}�;|L)�@�Vr�cK�����i�κ�n��ە����d<���=e�K�%��W�W�5QL�=u`C����tw��ӊ��l%kM]�z&I���c b���\���N�pـ#�!�D�	��/�t����#*Ũ�r}*��ZRu����^[��{��Ł�쑗w�+��vY&�b/�E�(	F�
�w�~�7Z�7����+^?�>l&� M���~���`����T`F~R��9�*�
�غu��4�(^	L8xЧOX��}����p��#��l�fi�<-,�E~_k�aL\�G �r����'Tc �裴��.�ڥ�,�s�u�������w�,o���TeDKi5�?^F�����/S�������y�	R�eݫ�c�'��cMݿY��Vу��?'�~���}p�C!>��3�BL�s�+i�[�x��_���[}���M�z�{�~Z-.׍q��$4A^�Z�WϚ5��u�yU����{�~�½�����Q�trS��|_�Ŧu����g��c	��6�K�*����.�ѬK
�ų9T�27|���#Ss;n�D�=QFީ3��O�	�x>*�J��VWfbL3銒�wkoH}�DT��
�k�W)�Y�C��bL�hL`W�N�Y��njqH3��7.)�օ�e-S�Y�.;�a�XL 	N�9����$���~h��1;�����8T�f��i3D�H�-XE��:��L�^�[J4�$�%���fdU���Vv
��V������ZDJ�~��A����俥m��x�u9�Ő���)ć��p�&]�~C�	ȣpV��l�-��d�����pa7Jf�=iC��!.�Efb�V��O�_e��쿰4k�νb��ᖒ��:�N�S���o[�i4�jo���Gk�C�m^�,��	j~�x�d���v��Qt��hH�չ��]N����Ɣ����-lanm�{�I; ��Hӭ��p1V9=��ن�k>��Qޡ4^����>�c}
��*�������7$��c�zS;#?�;��L4g�>�D�'�.-������� oT��1|D��.kO���a��/1�����A��w�g�tg�=����n�^u򬬤��^�I�C��Q�I�PU��#f�羨c9 !���U 3�K�G`�QWc��lTW�Ƹ ��n��3:��B�X_���O����:�j�p&,��${�l!� @��
��mEw�Ug��dQ��\T�ԟJ]_xEݱ<�س�ˆ)ۧ�YR���R�8t5ȓ������:��UH�s�x [��-V
�	�&h�R/z������i�8���g�_�/�=�D���$�|;��2⛡����Ӹ�w�\&��`1w��<���7��=%��^L�=��a���긲�A�pqW�&"�=�ʮx�=����r��9�-���\rE[Ah^��Er�A��W�ޗ�	������3:�E���Q����MI�&0r_p}^w�ä�����*�~$~�����������ؗ�a����,N�����q�%���WJz��åsgl):�X�Ԧ�R��d��J-���2c��\p?����'��7#4�Ցb-��g�4���I)��Tos�u�x���Z�<�$z�j��Ę0���Eԩ���A+#����Z"]��#���b��SKʩ���豸�.��=N���)�n:�Mj�gVl�Rǎ)����Zl����ͱT��W�-�#.G��Aqa��\���^��,r6�ԆswV蹌��RŔ� �6ϱH�}E�à�Xa��N@�)�O��������><ї�e�ּ���ߕ9�}�T�Fs��Z��Z>�ɣ?ƅ��)�r��Tq����$���v/V�f��k��=k�L��|��@w�7���n�������z��b�
S�vJ6����aS���������ö��\��Y�����I!����(;�2�A����Pv����q�_�-5>,=�fY����qBO_��2s��gh��s4�^��N�������bR����r�8��ԡw\ѰUiF���� *���G23����?�%z��qf�w,����cȹYE��#��$�򱴬x��H�]�_�\��Ҩ2�^��(N3)P�p���@I���fv�f�hEP��� ?0e�ǓF��'����}�� p	��-]�C{��/QjqLHt���CT����S��s6V�I����-���$@MrS���ϸ��ԥ��@%�~lN��\P�|jN�P�;���`��zB�� M.��;�ҕa#Յzh�sLb�b�ԅ�Z��B��)Q��Zd�6J����J�df����a���qN�]���9ʓ9�!��
�l��S�Q����2����n�_�8���e5+W,Vn@]*s��`�Z����ۛ�i�4�t�VH�!���n�}g�l
6V��>��8�g��A���Ϡ"��9�#|��>e��j�8`�^$Ӭ�w�wh|���I��%���1��Ȋۆ��ʪ������Hssm���M��^�"�8;���hڞ��ۂA{��5T+W��s$;Љ�-��|��>�w���C.��"{z�i�v��HC%����'{�?�C��6',)�1��gJڝ�O�F>K#`dkx���Q�2l�aT��}�� ����� W9�m%�+͗�`F�.b)	mG�%��P��i�iax`H�`��{�
jm�Q�)0��k��y����c���5����D�8�&f'�r��2j ������p�hH���Y.�����I���h�y]�}��|�QMH94����"3����*�[�����a<�_W6w�ٕ=aL��e��l������o���5�DB�}���xo2@X��c�e�Ϻ�����K�Q}�;��s�ۚIHd���J$$�D@��.�2�^*���]i�ק�yuI�Y?YD�*�"��+���34^I�ָ_��h��=^!)"v�#��뻦��=P��5�O7�O��
ĭ��W�l]��-O�:9�~���w�ͨ%���=�E�Q�~G�9��VS�6�v6���9K~��T)#|��y�������@D��S�kB?d������n��`�2�?P����"NY"�v����ou�=u��m�����P�a���æ�����҃�)����@�T�T�+����9OUn^U�'aX[�Hޣ����y��������V�^�<���X����G㈭�H_=�B�6GQ�V
a��?���m)��Wed<��
ū�1tO�!w���5X���ۓaGN�j��k���8�L�$�L�h$��WԔ���C8K|q4�n8�����E�x�T���:��ޮ���fX�َ��R�����T�����[.�T)c����C����'��z���;� ����5�N���)��\�j��8y�%\|hlVl��0��t.HaA�A7a˷��oȯ��~z�%	b���g��6%/��S�Nʮ�B�ͭ輔�����l{��E@�����K�"5��m'N��5�xP�[] ����[�dϗ�e��o\[7��~<r������#�Oz�Cp��#���!�`�G��چ��䫷��s����¢٩����mAO��mw�2�e��|�0_`�BE��3z�@���m��������8�U�t�	q8b�;���M��c���֦:���c\c9�V�j�ѲY�}�f��D=�e�P;�cᑽrZ�ml��L(ji������Bi;�:�Gk'�J��F�s�ԭ��O��bnW�%����(�Z���&��$}C�=L�%)
�.^v���2$�
����<l9��H���q&��������'0��%�ѻy� ��3Q��%�T�o��n0���L����)9Kt�q�`�%��J�}��V͉�����@<k�b�t,å^6��L6U�d���mV� �����]�_�'R��b,cDXN�C֜c��ܕ�}�<^$��T�i�����9AN��}�B+"�rk�i"g�¦c���XlxVHYEB    fa00     cf0�I��,SB������`Wi휽�t�LHXU��c}��0	*��)Z..�n���q�������ɍ{M�����c��a"!��}&�йBq[k+!۱�F�h�"�G����~P/��o��0Y�&1�,�_�X��4�E2Di�o��)�|q�V���%�sB�
���4IVs�iy��Ԉ3ǈa�W~[�>���1�ܛ<���@06:h���T�蹭kE��Q��P�H3x�?IW`b8d~9q�F<�CXj�XW��&��H[��.�'U��˗�2�����w�O$��=,����j��e��^���[����}���;~ۼ�>����ޔ#��e%�J�xq	�����F�;t����a�MJ3b��N��XLi��A�De�`њ�&��9T[�$ط�ܣ J���p62./��K�_�@�������ONey��&�S]����I�7��ّ���a�>B�D��8��#X8�}����cH�I�NȈW��ٝ�ȶಹyi�y��f/�)#���#�ln�ٓtKŮ_�]c�(: �7�,���&�~���=�I&�\��I~;��R_����<o��i:nP�eG�G�N���l5��êApXZ���g� qAÅ�W��B�d���%׌��fӅt�D�t�۱T7��;��+�u��nϻT�Cr(��v��&\4ߘ^���Xy��qU�4+�����3FIj_���S/�k�����CN�Hwl�)��юtf^�%U��aؽ���W�*V8O�@i���	1kt$�w%�|8q.�n�����̦8���e4�u>�J�/�?�5�؁==,��\�D!D}@�.jxY��Pv��H&�KA����&�q\���wC'4T��|J�]y9��t��~6��+e�3����78���Mp���mË+]g����?,>��L��1� |@��Cq�Å�(���6��/���3�>a��+���3�éX���g�K����YJt�G�^G*��ϛ�>l�O"�*I�9K�8*c@|]�صo҉��K"~��]�����
�U{�Hؒz����m;Tn�"W��=RXش��ݧ�M�HA���P�O�����r\w��<}g���[���\v���Z�D\��F�c�AR��b�< Uud>71"��oO���Ф��V(	���4rvD��h藂����[�O�������>h\�P(��y�FԜ(ׯ�o�dr�(-{�>%��+�$��y��/!D+N>�:���o򽉒��<�eO@\�k.��5
d�S�u��q���,�W/����w:�'�M��M���^��`+�@	���JKn+�n���I�zq���JΒ�TҮh� �Q�
L�xW��Q0�zG�-��|W4$�{d t���� �;g~��w}���I�O������+YO�����+����'�)fVW-LW �ͅ��9�
j{ރ�'�=�!_�`���O����Q"v����l?@�*mS������&�g��׋���K�`����;���V�$rh%�l�}�
�*��P��T=���f8��Os=���V��]Z?�x�����4���L���9�D���^��v��y���u� ɘe<��n�z�Jar"�S8�ȶ�ܬ0���^��#��Աpm�n��K��{��8���zM�4�?'^?�z��,�!�k�$7�Nq�z��1��h������N~�4���+� �~�FԪ
����e�P����<�п�lMj�@�X�q�!��{Ju�גʅQL:f��)�� ��<B�&�������;�Z�$O��j�Bv�U�?�0/h�;K�J���Բ��c�̡��X4�C1�b�A9D���:[�#-�y'6/>S�嘚�,S~��.u����'��?�'�S� ۋT~����R����]Qb"�7�����:p�ΰ9M�B��GF�*�TXa��o�r�a�Т�v����k��`�����?��ߔ^��x��kg:FS�7(��f���>�W�d��{�tFqF'@p���}�,`���#tԲ�K�0w+�!�A,�`T�(���,^�g�d�6��5�Y��C��qk�9&5���tyjN(�k�_�a�?���aИa�vD_�7^������������q<���/���|�JU��;��xC*�4k�;��-��	.,TK��UT��f�G���ղD��c��o�L� ��yyW��rݭ �ǡMgu)^ߎ�g�]f��(�"���}X�,�&��t��1�ô,�~9��ul&yY�e<5#�^ ���z�
��R�^	#�LI��6dH,�JAaS�H	��#�pc��T����i�Q�.�t%�|�gK�Y�%Q��K{��J?��J���7�c���0\�9tzڽ���FIٓ�~����,H����� G&�~��w��eȫ�J�o�d�����ӟ���4��rxcK
�[;+.8�*�@�򬃼����{[����I`D�k����HNRs����Vyb���0Z�/!C�;Cs��bgz��v���TJA���=m���[E`�X�|`�b�C��}�U���[�mr�W/�C�;����^;�*Q�y��:��*�*8�ϸ�5c�T ��V��ջ%�5�@ ����Q%|����z�@ş���?�c\ ��̹�P�#0����H�n�4����r.���CʯN�;�kA$)=���Qci)��NH3�~�G��ֆd�+���m�X��k@R�:{CLj^�zFJ��x鄬r:6��Έ�"\��R[�$l�࿨��8c3_�2Q�� F'5���Yj�K��=�hq�T-{Įu(���O�zun�T��@��\eh���Y�H��K��=�*#R^5_���;5�f�gA\&���f�]��?q��\B<I�	��@���i?��=~�~t�fi�lf��U̖E}���cY��}�qqJ�Fv	�3UT��#JD�/��%Y2�3���P.�ð���~��{�=�f\<4 :�zZX��2��\Xqgg�c���r	>O[�[�Sʬ'A#g��OL����Ŭ�s`��e�U_"څH+Bv�z%,�gB�TyY\�(؋��=�t:��7IȾ֝�w"����tަ��~�|X ��!ڋߚ��O�d
oQx3F3 !kW��4��7a�U�'�����T��/
3�G�q(���x��3�IJ��>���&�W�b�&S��٢�ʝ3ǜ��3�5��#�9!Ĭ��1��`��K�����ͣ?�i��ոT�/�mp ��yR�r_n�AQ'[x�Ĭ�+�{(��&#�)4l�XlxVHYEB    3981     4d0a@;���_~��bj�G}
����Y��>�ۛ�/1�Y�|�'���c���+��Ѣ�� f�`{G���ɬ���lI�]���E��k�ȴ1\(f���U���yx[f��!7W����6S�7�6�l�⍋~��?�s@ϰ�c���ǹhJ�#� ��.�CЌj�����,��LqnqZ<��V��3����^����$}���FtK6,�7���+��<�p�4ƴ��=C]�f`�H�+:}?yo��.vF��|��$�oq�O���h�珍�f��n{XGxn.�g#lReQ�;N;�����<�qH�\����,_E�RY�*i%�G
�̖}@��|�/��s��
Ѯ.� /���\���:�A�0����J���&�}b�8��꧞�ȓв���=n�cM2�~W��Xһ�&�\��+U�sR�|�?@~E�x[ef���zU�$�����mq�r�T+���*I��r�au1�MX0}k��"%=j�u6�D:�����F�ß�?���J���L����9�{�o(>����k��C��V&���/��Pq�2��Ɯ��m��Nտ�:D�&i�^���>)�#{�x��3�;���.����*?+�*?A��|H����Hw��Y����ZF������C���2$l!"C5{����&����j�Z�)�Э��R��B�9��k��UySH����aW�~�o�b݃J���UQ�j��9� �C�4Hp��C,*s2�O51?*��" ��q�.砾�M�� �]��DWM��6�uW��"ϛkt���O�����4�Q�.ʬl�>�p8�wy���B
��^�}�R�{�w�^<XI� ���Y�"��R�9�MR�����1��)n7����'��o��d>����I�COJ
.�G��ug�����ٵC����((S������m��rƦ`,u�gާ[9_gp��Q����1]�ʜHH�-=���e��k@�p"C��Iydx�s��;�6[+2����q�Pی�_���"�����~Oۈ��-�i���Z�k��%���r�.� 4⿕�z�CY#����2]X])�Zi*"��bb��N������%�D�eD,C�o��A+����2�j7����H�`RViK珏P�/�p7S���%O/�^���R	��Q��h��4:��,�>q|���&ϝs���)���{���