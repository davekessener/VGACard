XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^6/�Z�.� �Nȍ�#�i��A��A����|a*e����$��Cxϱ?�?5a��J@)������:���0nl��a���
�<U#��Z�E�d�o�h�7�V�?�G=�/K����nW��֛h�T2��!?O^��Z���^v�?+$���G��%�:&�㮓-s<�Up+W�K��\0�W�VH�����B�v�c�d�̄�f�A-�\b=���m}��8L>{qo��wO��
u�M؁ZX��x_�8�\x�F�6*�d�
V�u	�&p��V��F���;jOSl�į���<�]�A�VX�z�>,�K�_�Oi΄Գ�z���k{4�SM�+���H�F�mٴm4�M}7�
��I7�NB���I���ϒb�D�A�<�t3��U�E���mM�r�@�	yW5�f6��a{+�Zb�P�:l$d9iG�!%?�y�
Q�Ǉ������.�ਗ�ɒ�ܜ���Sd�M��,[K|��;[�������r����v
�^7�{��{�r���1A�&��8.i��ش�MR,����I���dc%��@ߋ�Y�?{��"&��{��T�r�q�nJ.��K
���J�7�,}�� cc[�C��X/0x��5�om!Qx���{ҹ<C-���Jg=��V ��I�j�ӌp;�����g���}#b��@U�sq����Ħ�� :����Bu�q��d^�7ū�j�Α�S������ΐ-[��:�D�n�ã֊�Jd��.����!XlxVHYEB    3504     cb0���8Y�>���"
Q�\j�(k4�i��˥�/���V磃h#��l�j�c����%4��'4�h��1|�;��2��S����[S�@�n���g��%.V���e��%̉�d��'�Z�# X7��2�8�"F ��Uln�^~�jR������T�c���
��ݨ���
\��Ss����fL ��a�}�ErZ'�F�|�)�j��G>����0y�ĹĂf^4�>�oAJ������<:7�n��4�	��(ٞ�~&k�8Z�m>�k)�>����|KG��?�r�ɑ�~'=d�v
-��[#�h�LN)�B��IA��ŚH0�56��OB8�Y��'���g�:<U�a52�J�ҔJhQ�S��0&�!F\�N���>���DC��K���>^��_刚�n��T���4�1�[|�L����h�t�6g,�O���@�]�r'F��I�f4O��蘒��"����g1@�k�-��)ds	�ۡb�I������T���\kg4V ��ŚG	G�|�Խ҉�)��4R6R�GcP4{��s�t8W��y{|���:)����Ԕ�Ⱦ�jS���	�	B�B��CK4!{y�b;��rlE��w�i��[��1/v���6L�G�����yb�s+?���e;H�\#Y�PՆ:��XC��<��ugS`��R��M����ҐJ��{E��#{z�������ۻO�L�c�4v�2LK�+�Pƒ�w&�D��	�����m]m��z��b�s��U1�k��6�i?���Z��8F<}Ļ^W�ʚa �����HX�!��M�h�f)D6Ql�h�p�dt-����XzXϬ❚�԰A	����wZ�59O����-y�e��b�,�Dw޸�7Ph2pi�KaW�(��epC3�4�Y5HO-ޡB݃��.	<��N P�bM�J5�m�7@��K礠��T�1���) �I�~$�g�|���j�>{m����(k�w��w��3\�5�&�_�}fiJy;�? \��ON��fX���v�D��h�'z�Rz�A�1�Vo�����x�t�l��E�B��,is�\����E.o��mRv�e8n֤�䩗�6I��[c�4�L�r_��"�^5b��H@����Q3�tLw���4��gQǖ&���Yv�z��Ou2��kM��G�9F_���}���h�����X�l /ig��+�����jun�>,_3\i�.�z�,�'X� ������
���@�v�8�Xݭ%������_<8���&q̘��f�()��{��'�U��6�H�-qv���X<��֜�:zz��S q)���I�!�$�������J���F��`+wŃ���H�-����qGx��P�����%A���5
� ���O��xoń���n�KSCt	=5߾N9c����V�]�;�U����i�@I�N�	������-Λ��Er�E�� \垌Q�TϹ߳L>�� ޙ�"(�sM�O�:��!� ��(�]�G�~��+���ۡ���M[$�h�}I ��̎(2��e�/��j�D�̱z�P��,Q����R?D-U�S�B���Υ���`���Ƭ/G�o�3�y�[����qW�}B�u�k��ꬣCy���d��k�u�C���c��w@'d�&ђ���!��t��PD�ZU!����Vi���#-�3]�^0X��w�<!�M/�n��K(2H��I��G1C����} �Q}[Y��6�6��j�����:9ӛ��\���A�\��Gq��m��U� _0�+��1�j�9���5\�u�Z��l5Z£xUL?�e��'���b�b��e6�*�dF)[��V>�O�+S��^�����A����D�SW��:���O��l���Kہ��\�����#�6'6��k���P�[e�x����u^_�"��/A�� ��w�9��dՖD�J=&]:$���5�����z�������:��o���������mݍ;��A6�*͏+����r�^8���ad� ��@���~�C�Ik��g�����Lc�j��=I�3V��T�uW
��g�뻽����-3&�B�`2	[mP	\���]{�5�T_�v|8[W�	�x�g,�|b&���!��V�����K�� ��#xE��ys���������o�K+V[s��1���Z:h��y�*u����6O�`-Dե�ߥZ;O����}7�;�Ut�"ҷ:��w��9e�X�ԅ
���M�� }�H��(ܬʞ�m�7�i�Z�t���p�P�s͞����D0)��=�3�s�w3��v��R��K�ϵ�r������B��H�,z����n��/�@)�#�6��/'�߸VViK�����~[�P�X�I��-�׫����"�B��ODq��{6�����HAV��{���(�}i��~,�DQ�#�yIF�|�����ZWJ(V��8��議ܹ*�	j���>���7^��T��8G]�.Ƒ�x&�US���!��~���֡%���aE5���A�C�/�Uވ�oϛ�A内sąRT<a��O�mK�F�Ƽt)s��"������&]���z�H�J��h��Z� im�G���M�H>��}�{�T_i17��2�#!gQ_��ax��Y�Y����[u0Sy,�n@�
������q��̣�o:��g!�g�	�Oi��
q ��ۘS���R�U&��P��`0�'r҇��;zO��;�JDm�Ȳ�K��{	^P��Hj�\mҮ��~�m7��g �J�C~)�Qk9e����Κ�������\��>�q���" sC��?�'�h_K��.�mT</˹ /7rd���Q�=���x�KqE��3D�HB�������.�t���c�>��b0d�CX=T,����d�������(��/�oa�k�������2��3k��'3*u�P���*G���"1[F"纶����Ro��<֤S��!��~\Q�^1�NU�������V�Q"i��T1�8��j��s�y'ޏ���ijC ,{�g�l��>��S���_�-Rm7���R������i���K�����U�I�HQQ��;�h���}-�Α|���l���o��5�=T�c T��4u��)q��m�8$�M�*�a����f{|}[[�)��� i����L?f/,ԐX���p-.