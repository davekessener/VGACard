XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<����̈́���3i�l�� �鵏�W�{~�i��|\+ݍom��L�q�'�gϐz�U GI�@�6�QõC�aS>�(���E}�>wUw����q�ܟQd�2��u��]�J`�?� nq��s��:��%�!Xl�v@?{�.]�tF�S7���f���#C���6cp��T9?3I���F�EhmT(�e���x��S�����L��,j���RДC������Mޒ�W邡A-�@/~I��AUA�����qB��XF��`�^��1ή�*R}���s�T���}keBX��{��x���2
��㩻�0z����G�Q���6q��PCZOA��a�4cT;��6"����4��P(�/
��,��[,��%����d�I ���;���Ey�����@[Sl�"�{�X�M����Y�p���ǆ,9���y�Ӄ�;B�&ӕ�CSZ`�/Di(�}Ej�	��Ї�1|c�+B��[�7�t@����Sg{9�gl���M���$�D�>�Vݙ�9fo�<^��R���n9C�?M���!2>��$�\�m��k�&�B�k�P�`7�?�Mw�T������F/t���]_��2�)*y�a��K@�I�����PN#2�����-���~c��<��~1��3��>v����ei<}9N)f:�����~83��iz44dܵ�!*/�mS-xnJߍ����d6ͽ^��ڪު$��.�m[�G:���|�B���f����X;nC�d���J��F���Bw�QXlxVHYEB    29da     af0o�֝�z^psfz&������S~<�lS����Ò�eC pv�'kdpD�*����|�*/4쓛�@�r&k���Q�c�>��4�#�F�6}�M ���5ӧ���I���jP�Lb����I����7u�$�<�Dz+�.#\Q��kP�JM��@���G�BOb��"�ù�-�	�
��c���)�<kOjʿ�3��հl��B	I��� ��!��[v~oF#�D2���W�H~�T{V\�o��z���>��\3�*��'ٺ8L:�
�<��+�����Ӯ�2��W���)XCzu`ܤ�_�U����arJa@��}��l�(Y*i��4*{��^ފr�?A����c��)n8�G�}�N,�GUI���pv�S��U��O]�~N�xw@t�NT�dGٓ�cǧ,������E|�mPy�d��d u�엧�~�1�|�x�yȸ������s� ��u_I U&#�$U)L��;�Bx�V�"���72�z��#�� W�u@}�{�G��_��S�q����'j���Bk%>�>��0�~۾�T�VVxZ
�.��������7�����\�a���d��S�^΄h�Bk��sݢ�l��N����D���%�nA�;s��:��/ues�:ea� ?��}k騔�rP��c��ef8�"�
FR�O�V��#�{~�`>SD�T��z��T��(�4Q���� '����	q��f�@E�?V*�Y��@5���[��D$B�Ml6����3��Q�R����$ P�O������)>k�[�3���1�6���k��p����?�1��[��Zw1�}��G�- Äd@JQP���\{�ي��3�O�1�l���<��`��,���S�m��T�V�xm8G_d��!�������W�:�7�B�K���*�8+|Giϝke���A�S�Pt��Ó���[�`��*���U��z>p�!�s�Х�K�LqC��*EAP����9�O
(��|�b9��U�$9�V?8���3�d79��)SN
�'�cȽ�TS�<�4Ӝ�FF��"��N29��� ���s�/�y\F%V4�W'(�9�:�H���neQf�
|`���_K� ��� ��o}�d��1�%=�YW�b�����(f�ͥZk�.VR��#�6J�Qr�=��>�g��a:+�K攺�G�0*�چg�����ga?ڮ��S�P5U�]��$��m��Z,�%���j�����~AF�8��X�K?7M�F��qx��N������!)����;ʾ֚J��^�/��zt���Fe���ռa��z�?+X� �C�A2HF���bT��A��g�ñj�-c���I�!���# *�8�ɻ9�{TX݈���d���Z�.�P�o�F�=�2�]�i��cIo�,� 	����	�g��'vU��z��:�jK���B ڱkM��/g�u$��vO٦�~�)��\_QB@s�ܨ �x��)j3��W�}c<UvM��AJԬ cf�#��"/����R<�5y����?Q^2f�u��}w���jo�a��L��P?%�����)�\��-'m�W�lDW�*��քA��j�"����Rp�Xzh%K_r��sW��qr6�>�K�}�@�`�z��Ϳ*_���N��Zio��i��=?�c�`���a�R���lU�K�w�w���m���RZ��9n�p��	�G��q�bq����Q�u�g��A�S���ƪ�	ĹC�H�ԬE�c�\f/���ڂo">��a*?�_O�����'S_�ڦ�y�-����C�r��B �F��9my�O�UU���AţkG�e�Ag��=�luz�o�xƃ��:٨��`j�qR��+[��'Y��î�eA���B���MϬ��sJ���y�&�tj>�&]x$���c��L�"ߤ��\�9��ࢂ��}�0�Ȭ�i_��7hGb2X�T�V�ZKk��g�c�\C�ڦx����U[��u��&�DT:��SnMO�T5�r�eBr�4���'�&|֫���X4����N����\�V�ʎ!6�mAI�.$��ҮԺmmJޓF��[�:󀠵����Ys��ʳ��Δ����Z��;a�e�aN��8���V?^9�Ć؃�w�)!�3���C+�Sա�����}FMꓫ �B'$����PB�X��݇��^TVI�xہ�����z��+��\���(�Uh���]��W��^��֪	+q��o�ӣ9
��|�$$,���0���W��T���2Mu�I>}f�w�`�I��tM}~π���e`�Y�6K�?��R���ne m���oVJ�^s��ƣ�I��\E������)����2҉���ĭ��"��q{�*~"!Ea�B�h�1@FL��m*)���z!�'*�<�F����{���F.����]�bÕ[~�X�7�yS�! Eb�͕���W���,T)M���!.���A%�7
�1JX�WU�\�1�SH�k8l/\Ǵj�l�v|q,"(�ŵ��=���R��9Z�ئ��LNk ������зJ�@�����35J6p��Fq�R����r-��t(�Q�gTʆDk݄п��<47�*�������4�����GT��"F�������+�ܖz���M�3%�&�/z�2��J�ӆ6[�~���}�7�Z��n�K)�n����/a�����\.׈�"���դ�4�P�2ڠ�+��8��ZWe��L�䧲)�Mo�6P!��k_kZ�Fs��g�`��