XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���̸,Ϛ�L��H�U�(�!�v,�Xa���&#�2|��\3�|�}5�����*��A^#lav;|����EK�B�d�~L*sZ��9ƞ�5�w�V��?u���Hi(C-����9��\�Ab��<H�i��!Е�e�,� Y��J=��c���� ?ؘga�1I�T��Kۢ]�
g;�WܴѼ<j���qMh<���Hs1%,ތA^�ګTy��-�_�_�(�Y7�� �B}�I�����v���IZ|�g�	���9��٠��n ,?��:��Z,N�A�0���hQ.��N�-r�Әb^i;��"�(b�>���[}�RX��W�\G��S�8D�\�'(�>�� �����`n��a�(�H+�<}��;�(�6�����X�n�q�|�T��G3�L��{�����e�f���0�K�-�Goi_,���2�t�0�)�\u�{�~��� �K.A��Zq3u0��\�i�)�^���r{�I�����9��#*�<��9�?Cj��ባ�q��;��m�kb!�)�b�!{R�'��_[�7���Ǳ��XW����� �С�{��6�U+������l�\��X	W��E�N�.�z��ra��y˾i�'e�ʦ6��M+ R��e^�8�V��dR:
����Tq��� n�>��|�ps�ۼD�f����V���]�bm;^dR$��Pl_�Ѳ:��U�(��_y��z;(#
��"�=�jx�5k+ί�E�<�C��H2�5�%��<�+XlxVHYEB    fa00    2480̈b�j�J��*��L������+���%��K�L�j1RG,Q�/��>>�?c7��k[�]%��@�3/�W3��z0���L�
��ZK=�7��Q�������`?ύ��]V6o���H�-`њi@���P�;�=[������2L��nUQ#����������C��w���T��<V��H�� F��.��Ȓo=m?����ע��Ƨ=;�C�?p�w��c�E�5+���o�8��+�0LZ��U�Y�����h����k��;����N�Ŧ7k��(2�.���g5�~���'��1���{�� 1����L�����ǥn&~�A��(�D�ǍY�EԿw�� }���܀���+���������?+G��ء�pZ|���-ĩ��o/L6|���,���)�Ө�5�y�1����ά���)ql�{���%\���r�8!�+�HDX�E>#񰀽�<+��b�\oHP����^���u�U@(��Sw�0����j41�ҹ�v�{&���\���?XU���=���Rx�^X��z��>T��R��=��3�3�.3�`�x��%z�;�<�,N�vI�I�$$���ᠤ^���U�Ȅ��p�#g�zJ-�΃"�40fJ���@���C��\ܐ۳��,��[,Awra�bA~���~�c�������/�m@������f����S��*9���CT`E����}C�?aDZ]�E-"�f�-O0(�~��H9�D1�Z��(�{��vy��U�Ý\5ʺ*���̳a+�����|Ժ�x}4NG7bO��ZY���s��ij+�n����R"˃�v0B̮D��*��}��=��Q�{�����*<*�7bZn4��F�zWV��v�8��%�jؠr9U��&bi�$�<o�ɖoo>	�
�u�s��8M,BkV�ƛ��3Jf���\ى.B��!�xC�3N�M���;������s^ ����zIlӍ�-��r"oT[�6���^#���D��HV��}k+ق=9^��.`}Ns��r�9�٪�QJ���W^�k����w��bm�b��#��@�8�E"�&63��d�h�{�=ݡ�3߀�5�`�1J���k�J:� �(3ܤ8�n.��w�0�+����I �+�h��[`����`�;|9&"=F[t�+��]�1�� �����^��ܤ���6�ĩ���1�u���B�!�@��l�r�F1/͟)0D_ZJ�J4���?+��l,<��#��{8�7����_�������a�hCV�4���t�4�ގ�{�80�b8�O��+�*'K�[��x�[�X��^ӡf4��Ui'�/�4|ؠ$X����E9���.��R%�:�(�������2,컎ڢVD�c?��G��F��S&:�7ΒŻ�`�q�%^X�{m�ϵţѴ��ۿ~���C
�N���)�kz�r{L��%�ʚ+���H�lcٕ�mn������<����{�t�&v7/��J��/��K�V&�n����.�^��{iQoA���Cpu#��M` �T�Z���'9��-	��@
h/��x�F��ys筏�t�� ��&����9R��`�T�*��V>��u{+��W:R�5���O�Hn�\���!�j���,�z܋��2,wl��|��#���%�z݈�m.�P0��1������P캯cS�On^���B(��9O:<�ADW��m��D�]z��$��%�lm>���[�T���$�����Կy=wfo�m)ᢳ�|���HS��W�)ƤY�f|]����G�	l���ùA�P�0���	�A���q��Iw.��o@_o�LIL@[ژJ���Z���t���.:[�H��O�~���v��+��@���@-`��Q�\�2��x�E:Q�iu 5�t�F��F�*|�L��P�O.~A�SC,q�#`��I�=}�qɃ������g;/}�+��B�V�`-lt��+����I��S-�kp�gCR���W���Y�ߊ8���x*NQث{�j�mS�((P�Ps���]P)W8�cק�j�
��� DJC-�=���a�àD�+r|��ٮ��Vv�(�ᶘ�`j�
�5�y���%�����@}��2�$�Pv8�!��?�gB�ԃW����rt�E�.����&^5�����3}��`�G��?�B՝ISAͮ���<Knxӣ�$'�쌚�M�Qn�E��a�n�+��Esu0x��5��u�"���(K�`��N��ۀW	k#�-f���4�[��?��
p����Ӣ��r<��}�o5K��h�?!J��Z.�}�/r,���e��n�҇��_��f�Vu���ν���a8�f�!n1��4��Y<�e���A�<���i(8#������I�q�h�3S���<s/������~J�>�Ju
ׯ9i_t�}�'����Wߨ|�j4F�(�4��?Dl��ܢ豔s�Z#`ˠEz��14����j��%��:�A�v����^�g�Q�Q��v�!}j���-C����`�P�4,rǂ_3���f�bk�X�.����]Ch�@i7���.g|��*�[t�꟝����s�޽���K�K�j��'}��s%�N�I�ҽ@��wtQ�C���O7�v[be~>gB��2�� ��¬V���t��(c���UC27���W��X��ڹ�����48~�8_���SC���r��n��Sk�u0A�����|�����.�#E%�(v�La6m�5��e�N1Ф�5��s7�m1YK�y��~���
n��W�~�!��0�N��[VM&:�'�"gV�?���q�*@��判���ӣT48�^�I$���%e��W;#)#��9&��ν�x&��v0yEI��z�u�f�U+��[�7Dy�<��;������i�E�2�b�*� h$r:h��ϩq#���zm3r�y��*��{�x)@,d|�dĢ)����i�;���y���S�y����<�p{
o��R�v?<لF�iK�(^o��F��?��,��=0�桂Z�d"t5��|�1���&nc�1�;� �lY+������>b��C������[�.j��9��9��y;6N�:%ǋG�HSPFjIFqm�GsJ�<�w��͋�r� ��8�M����Bz���ވ5*>��\�>���)�#N.���ha��J��7NTK�Wޢx�)lzp��tζ,܉N����ns�#��F=�6�CPƢb&O����({X�vq:%7E�w��ŗ��1i#��)��NS�j@�;���v	�[��j��b|�ݥ��A2!�~f�6�R��5��?���}fG��և�
��@y<�����>����1��$n'e|�&3���>x�������H9�g*+�T(?e�u3��K�)�6+�[����{_�v܄@V�E���T���/J��c5�v2"�}}���s*�.��g�8&�9�f����i��ٵv�����YS��.w�(���v��Y��k7=�y���-)�-gt��WlU���4�4]�i���i��+�eF����а�x����x�	���n����M���=����a�,]�tC4�_I")_^��ʩ��G��OeМ����h�2;Ʋ~�scw'�rh|����%ܿ8������]�ū@�h֧�:����p$i�I��T��YE8|}�n��`-eD�/{��k�	��{D:t�jV���0}d����{0���F��,�Y�WN)Z%����^2�.a���W7�f�P�VM�;Ȉu��"-����E;���r�3�H�2�::Ij�*�!�Kh��ޯv����?��^�;}���>��&:�]��
�F1+��|����:mN8�����)�t�Z֩[���^�z�'蓳��!�[9�V��c"��_1Z��]�����dgy#�f/��}>v]�w8Yz{����Vn��c-ح *��V��o  �w�e�m��J\��o���n�X�"�&�N���Q����m��T�g�A���!u��>��ʌO���=�,�l���CVL��d�O��8Z��c�$���\�)w�}��Sz`��od18��~xK�!nH�4Y���f]m�/[^Mɪv4m��[|+�8܊J&����oP�IdKB
">��|����ٲ��7��Zޚt��Mv`����ύn�^�9&��
� ����<���hl�����p��ԯ�0�-Ս�{�cx�E-, �Q'�HD}�m�������_�� 8;L�ME���S�Zom&bzm7W��ۙ>u��ME6��E����J�ݐ��}I`��W9�D]��	O`��FW�4��{'e6F�
��g�q����a��[~��]���#�y;K�<�`a۠y�e?鿜\��M�c������Yr���$��mf�z$�m(@3��	����5���_c�Q�R���ܷ`Z2a<4n���B�Y%���p�����3y�	�������%�\U!��U~���Ѹ-�/�OF_*.A�����׫d������`�=G��i������.�c86��j��<�!���H�c���]ޢT�}����J��rJ65���F��ʷ����.����a��k�C�19�)�l����p�)d�.���g;�6|�H��~~�Kht����X�e="w5C/;W���h�e�����.<�����^�:�+�2~��@�2�����_�B���!9���CAGӷ���C�'bkx��Qߘ��|/.Qu�`�Uo�X' ��"�]�1�u�KB
��
�|�&�Agp�q�́������
5&�Ќa�&�RpZ�"e�m��f��Eo�ݡ����ě�x{�Jm���g�Ր-�?����B�\�Ƿ"Sի2����}�X�m��˴��W��5���*Wv��aKx�����5��i}��V�ɯq�3�UT�T�>�"�Ze˗i�����RaX �:��ۣ���,�D���l ,��`n�n���=�"���x� &��l*�p�y�A��.�x͍A�x����@��-6)�O���ѷ,�dc����_cixl�i���<����/�e �z{'^h5���c�wD���`���h�z̃1CI�(�C��nw�iid	�-�e|�@�eePZ��%�`8Yh��~�~[g'��W�1_�H_ ���
$ ��6`�zNλ��U[��s���K�\�����@�|��.�2��!�����ͣ���ƒ��'�g��b���J��]�#����UʾZ%m�b��aV�Z|��Z�/bA��� g��_��5��j��*h7�P��C#��7Ô��X�j��8D5��!��t! P�D|����e쿰�o�9/��D�a�^��Cg���c�����(�z� �X�
0�M�P��Y�
!���vZF�=�
ܢJx��؏��vh���P��n�@x3^x]Ϊ��QW)ښ�`X��?�Z�����l0½��c��?
�$���]A��1ȹ�|��6��a`�SãH��%�Q��$V@yh�>�pE������k�5�ssH ��'�(�+��z�)�<�F���7is���i]�c`΢&}���d�)y� ���og�	p��>L[�?jUXCV�,�L@/y
��[-�8�t�f�6�u�z�kY�����g�Rkq*Q�F�T:A��K�$YxDbO�ql^<�2�W2����G�z4�N8QU�I����>�#Hg��c�ˈ�z9��]��1�[�`�0K��^��v�O��")T�ۂ�(���!��0(�wn�Q�h&��f���G�?���:�:�eSW�Q�Y���X�x���z\\�w$�Z��s򉱐U���iO�~ �Q]�+J�}��F�}-
���kj���Iy��Z�fv/́
�!�Y�kv��^���|�VJb�ԆP�\��:l ����Cea�D�e�aH�	���$�%�*�tcd�9�oOb,�,8���ƻ�7�7W���-+0/@wU�8��D��95Gz�=r�*!o{��|�~[�oǖ?#���C�h�b�:=�ê�Ʋ��FWL_����R靤�%ec:R�AQi��y� r<��-d�N=�tA�`F��7};�s�Ӈ�ͷ�sth^2?�����U`�:�8y8�락O�:�Pٱ���݈/��Q?%�a�����5��;�9s�K��������΢Ǖ�g9K s��-���$�B�ݳ��e�6b�3���e�U�u	���������E.�Ns&�~�O
N��c��;Eߠw�Wނ�~�c�z�ԡm��#�%0�e��E���i��!��d2�5B�J��x�k6ܔn͋�ЭgfE&�8����A�f�hx�"ȳ���I�*��Z�m��7.���e\�B���IǾ{0���Է������[4/N2���[���|�� �Ϳ����?QbdN�B�T�B�����`3��j+֟O/�Ʀd��|L
/�D�*�.c夹�����P����=잯ˡ
�Xԝ?=7R[���68?@�a��ZR���_�S�i$�i���m?V<��H6����+r����-��8h|}��j8���%���z��A�Т%��_�n��cY��f�<ޭ�;�+�50zMI�����
Ft�A[���<�Km���o���R��g�vmvJe�[T��moRN��.�oGW��1o�~[���&Ȉ@��V�$|��8�$���!��إ��Mlw5���He�`HHe��ʓ}����%�۫qR��X�s�y��[�
��Q�D/{��:zA:�,�'4�i�+@�ET�?6YK�{�W�[��'���TB�6�n�L8�w��̽xd�&{�Ss�N7�7�P-_x��	��H��ecӑ�Yg�-^�}m��I�]'��a��<�;x�`k�L/�`�����l/]N�v���g�.�}� f��<_�25�#�#�"�msh��Z���m��$3u"Xw�	wN#����{�� �Ϸ�?��7=���T�����[(�a���E��5�|��H�����Mբ4w�dV�v�:$�>��iA��#P��] �T���	��y��G:E�
�qTk���h�b��|) O������ �T��u����X�5]E]�V��c�(N����ozdJ���m:/��H�����H���e~�0#72t���J�G�a�8�?�6hjݗ4v�=?�I�_XZl�D]N8g2�-|V�}5�*HL�ځ��� ����`����!��݌�w�������djQ)��Q�2Ԍ2�"|ֻZi���ϒoJI�}aл�H�]h��ڄ�-��<�,��͠��^��뙥��	�楡@h�]>��S$��
��N��$�`�%X�Ó#�/��zW�x�jª�3�ϲ{���@Qӗ�O�K�P��=�[�4��v ���Oyy�2IsD��Үvn�(��*>u������:�B���;k��ɨLԡ� �f���O�D�u�4�xh�Cgl�s %'���;8Կ}1x= ��?���f&6�U[�v���la��k�S 󡜇]�BjeЮ�\"�K�����v������èFe�鴡���$ׯv�}�>q�]��2;�^t.�p�Q$6�R�`���H�m�^*���4 �Yx�l9e���y1A�\�nɮ��<N ~�1|n�C�^�I�N��b����M����\��z3��f�)p
�~�M��	)�"�`��VL��.�G������:o��L�N��\��6R���_�CVz%N�:������,��/��EPNе8��|��Vk���Uo�F���]tr�jۅF����$پ���@�)Aݖ��gm��U�m���b�҈���#�v����q��ӿ�5�R��t~�k���ist9N�h1+�uLN%�3t��8z�7��V�y�?�G��3�j����I��8qV��C���]X^K��J���7�Ʋ�r����r2�s�i(\�� k���C0���/��̷<r'V�sg�T"� ��%�'��}��
(�ympX	�����w�	-O�eoj<Ł�̛8���+���TO8��K6 �?��Nܼ�ׄ������j�j��S@A�'Vs����:�d�����r#�В2��	�o��."UvT|�߫g�|wb%uSi��A9�+�8yJ������XJ����b��;����/Wg]���E�8��#�;X��l`	�0��+�n�qL�u��#��6q��s���L2�آ\J�H'���3���5� �;T�^.��z�9�(��$?���c���/��̞q�{�QM*��3G�\�����/A0g�;�yޚLI���@]CFl��NW�o'e_ǽ��I�湆`��i�%-�2t�| 3����|e���b׀Wob��G������Nnu{��3[fj�ܢbl��2�i������摱nӽr�R6����������D�`�4�.�Y8Fn3�c}��5�~sb�
��"o��-�)�F�:�[f`�����	���FK�{̶��f��Dh�-���c���i�_+#�L�-���z� �^R�q�`�L���� �j�	�2�?:,���!�&5�:9�7
{MǗK�JR��BhB�ͪ�;�Sp�	8���N@�8�b����A��^n�mpkT�_/?r�"5��'��������Uu�՜F�c4�^�|�i^̑QcN����2Qs��H��'����������������������!�Ia�+d��Q[�$��Y�I)d�K��y�}�E��L�6�$A_���z��˷�Y܈]�_{��:�j���ZHN,�V|P���`���F3 -. !9�����yZK?�x*�FyƐ�~`�PP��MBݢ��SN��]H!���d��}ۻ�ֻxGy�2�t@��KK֤,�f�&8#M�J��W��]�����m��*:��b%��\�kL�	�D����iy �y�z0)��?{����,��T��P�Wlw�wPz�T��f���<�u(C��{v���1��LX����a蠀a�.�k�;���e�7^U/�����ԘAY^A�:�Vo���=�cxq�\S/�b�s��jJ��~�]��M�g��-�����{��t%���q� �p�O�/��Ŏ�#&�p��%��B�>�'�u�6�'yF�M(�lV�WE�9�"�����B0�Q].�l�ެ�XlxVHYEB    964e    1150N�[�Oh�T{}�U�������������;ԅ�  ����)?�k]��)�$����Ť^�PB�iGp8�+ +�Oŧz@.�N&/ߖّ�J<L���k��x/9�ΛCv}�`��y(˒w�%xK�Ma��DҊS��T������y�p�v�SOax�(��9O���Dgd���Y�"������/F��s��#�+�~W��)[� cי}�:F�F|Ň9��~_��Δ��5�(�0�yPف}pӓG���h��͟�Q��B��8"��b���`�<����UjG����y;��! .��ڈ��yt�8Eږ��Eď{���8���pj�c��͊4[�e����2h݌C吅�N�kɿv��Vq^`&X���h��~����u��j���'Ì���#�3S����1eڳ�rͼ���V�аn9����դh@e_K�v#����9Τ�e��<�d�ٺ�3�s��"CK7}�&�	÷��j��6�Y�K���C��1��%�"�Xmk1	�E�nd�vj~燽 '�<�� .�n�CI�/����;��*��)2Lm{�ށ��Fy��왯���!q0�@���t�``
!t��Y���Q��>� z�m�vt�f�9��k�-�Ɇ����ܓua��D�Z�mb<�'��Y�Wb�8���S0��~��|� d���P~v��:9U��@ڗ;	�h��e�����^%�# 5��n�<9e�$J�%p�)#R	F��C�7���2UeI���Z��ߎZ|�>I��aRW�a@��� Ƨ�|���=<�I���~��_��㱦�0\��\w?�q�I�\�,�]y>�ltq;+>�7�{�K�m���8A�L8����I��L�8�1D�D����\�f���*�#��Yk^T�(���Wg[���A��A�� ��fE���c#Sڬ����%e���>��T�T�e@,�l�LYէW�w=���YQ[�9��9�!�̃ݮ��
5/jJ�r��.��}WHf�n��~t�<f�!��;���$����m��-8��b	eѻc�F��%���*��������%����4�u�� �����%�v@�߹J��W���J �'\�+P�l��z���mP�;�4�RӴ���C�֯���ʟm���\�xJ�1�#��j�YPq���ri���o��}⣶X��E�aBz�nзDC�WQf�9��Ƕ��J�H���%Q�0�ȕ��dʿ,]��A�Z��qbУ5�j�K��#XM㓍��{:��z�h�B�#KW�)}���^��|Գ}9��+��#���rP
a�69�o�.��Ϙ�d������Ed:~�[�q9�?,��6R�D1"ဌ6�X՞�ҁE��������oK�[^�_��<ZJ��*�"��.�t�(Aqȱ��+r�S�*J�����?aK���&��In�2��6q+�!��(w���VN|y�cY��A]Hm�ގY����=���I�1V �z\����c �}J|�,UV͙�~�ǲ����Ӵ`���<Z�i�iKC���<���G�u���oo�R��;�%���"G�s��9�����GM�Ur�u}�ST%�2y	W�*|����}( 0dyw�͛"8�i?�g9Aq�s;P�
!s6<��gm����[Qo�u;���`曢+S/ꦔy�=.t�"�J���Sɾ��	��BxEߨH�Ĩ��"�}8GPC(��k/K�NV=ϳl����G#q*f�m�;W����b1��\�pN���<h�G�O��l8�XF8�ƣ�Y���#k_�O��.�A�.!�/f��_���?8�$�3��^�Qr�)�L=�>a�vX���ؾ�)��w��5�a�c�Jmf^H{#�W��<<��.5vyPWӤ�����㿐o�D�+^��)�>h� 4�\���6������OM��q!"������'d%�t1@N4sa�wP��u�Y�ȇ8��?,p�!�F����-�/�fFW����M|S�����~�5�ƞ��vH���nh?ȵ/+�����M{Y�{�y.�b�q��Ӓ�����}���G���b>Qd����p(��>(���"�+���i�l�U4�f�d��HB�X �����EBT����OD)&�6g|�
gN���k@��L�:}�"��gd9�}a#�U�b��yr�񴞆sd(D���6�������[u����U�~<��F�t��yd$��e��=z,b�`��.�ʑ!�}�:��9��7�+�SOt��
Zn�ټB���t���A���[�蕗��P���qt:!~���@0V�H�*���t=�f����~�P	�ij����ۺps!�gʏ��v7;�XD�y��T��cʓ��`I�AY�n���I�z��a���'���N�憕;�1J,����̃����ѫS�f0y�G~Sk��/��I)��&�@(\W*`�r��pX����0��J���3?<ټ��'�}+k^�5�ʣ�W�?d]�h�� ���sc���!�o��r�t��LϖGO��؋[A6����r\7�ݹ�P0�<��џ�}��pH��49��1�&p�B��z� J�$z�g����?�N����Ù2¹��C���N#�2�7m���s�@*~!>^=��7�v��&�^�&�eg��
D�g
�r��av�_61t�u�I�hG;Â�m_}	���u;���Z��M
����������HD��P(�fnŘ���r�愧G-�^��4.,����1]�y{W��y� �[!�:�M����_��w�̡��C�q�V���jp�<Go��x��7BOf�u�PcL�;Ȕ8@H�(�-%b��sP�u/�D���(�����I`8s� R��)L%�	t����|��r�V"=����`ʣc�G��>�?�P�͘�P[:�׹��+������]@Z�j��딱����ޓ�����@z�GB°KZ�"�ߺt�'���(ƋH9?bQ��@@�,U��-��K��g�nW��ce�[��Eʡ�8yN��3��аz��I����S7C>�U��<�K�������\���uu~��zZ9���V��4_����NQ��Q}ޱ,D�*^���x~(,���_=���]��Uf��4B�Q�P��z~�R�0l�pr�4���BE:�A*Wn�wN�ʤ���>��y���Gymu
U^��r��߲�]<0��"�S|��I_��3�I�M��ڋ&���{��}&���Ǿ*�S4����Vcd�c��6�B]z�#�Yj产OU���S&h��	Ot�P�*'IB��j��(d���??a��$$tB�I¡�X� �ek���Afak-�j��ɟ���b�V�rN�[n��c 1������a��K�r!��������:ʄė�<ev5�ꃤ� h��� J��9����+�*EP��8 ���'�����R
a��M���K���N�P1yRc��A��R�4��� �FhC���]:lJ�0��Ķ��SF�`�kh�@M�k����a �݂���bp���e���s^V�m�Z�@2�5\
>l)�<������'������V�>������^踂L�u�0�!�l��-�C�T@�O��?�
��ޛ��Yc^�Q�A?5U��ğޥ�(��4A�bh?pZ�-Z%���k�I���t��{|��Q�:��3v�����o���!�.���]~�'���+��iD�M���Z	�І�;�g�Pǐ�0��&���r2<C�*�bc*�L�}__�U�b�>ϟ00y:�D�G0i�(5��}JOyj���M]����|��R��~����sp�����v@f}���c��V���6��̠5aO5)�˥�QJ�x2I�׽S�cٖ�M�̭aѡ̅I>Ը����-��`��	Muy@�w'�#t_�E����q��3˭sYpmg�k	���<���N"���Е	ږ�X�*����o�&g��(Y)�oo@�Pw1��Gٯ"`l6a�%�Z�ɠ�C��3ql�0O�a��i��Ў	+��#�v���$�YB<:<#��"$>M5��9�y`'��/J;�yyT�HŚ0w�� �9ȌR�P�mg����
�K�t�T@�5�&����:�U�E�g0�n�����Xt! c���0J�J%˩�܊�#e۬]2C-r�Ȝ�1�T,��)4�d&e�V'�F��Ze��;:�o�R|sM0�����ύj|��8(ϻAx��E�TKW��s���t"f����\�{X<k̞�bZ'\�ȃ���yr�h����Ŭ������G�ِD�DTTw�})"�13Tf��-�TF��C�I�K��> �z��A��)U�FKO7��a��3@�j�j��yg�b�*�F