XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���,�qX�a�WU7c�VұA�m�oHj�Pu(�T,�����*)�7��/�J��<P���DS$8�I�7Ȃ\��Rq�1�����-��Z[΁}��,��I����?����p��b�+x�&�[�]�&����`�����dY=Z�5bk��mF�|s�5 BH�:d�B���a*�C� 混�t@��0,0!0,!%��ݺ����R[p���x���|���+'��_���_��v\�~�!.ns%ճ�ž���G��NY��l��-��m�y4��TFq��g�9%��Q���M��0U�ƫ��` �FL�ą������C���G���_!�2>�ϳ�].�'�?��]��)��Ea?�eP�h��h�g:t��$���5� Q�����rB^����s,�_uߚ}�� �S���H��&"���<T�uHJ�jF��j�?�Z--n"[�qu �?.f�U�,oaբ�D����W�^�*C�4�qA4�(|�5X4����<�,��:o� �d�PE~�^��d 9
	��&=�te�`����M�C,a]#��va��o�H��^�p���r �
���l�#��5ΘP\�a���H�z�`ۡ�E���9,���b���J� �u�����-���������AWR\Lgќ+D���K�7��JlA���[�Tu�HT��l��&�J9��� ��l3��'�D��Tw�}R����I���W�xF�ָw�����;l�?�s� rt�0�K�+PT��z�)��]_�R��?@�XlxVHYEB    162c     850�h�;q� 1L�ˇօh$t���m�.L���/��o{����H���gwqc�����,O�.$R�g�U�O�O��$��Ce�5
���(�#/E�0�5>��<���K@��U� o�g����&�>�c����z�ۯ�}�1z ���	Cz�N��E��>������9�����*Sh�C�5���兩E�����ן<|L�@n	J6��
B���tؕ������s�Ԕh�)m�v��O�|�H�#I/� A &��D�W�#���PHH������Hw0��,<��-K'J�D�}�.jߐb5m����5V�I꺍;�
}�k���!����p���4�&� ������C~.Z�R�K����uv>��\� �@Q�	���Q�a����j����"���"G ϊ�a��E��	��Z���E9ɿ2�w��e7|5��0���NL2���BN��EbQ?�c�I��_=Z|�D6�6R 
V�Xf�����I�:e�Uj��ΛΗ��)�0!9H�wC��\���R
�F}�9�|7�'Qjn�V�s94�1M�tX�jov��%�?���ߡ;|��E�sf�fa��q�(�|����̘�op���e4n�\�rp.^Ar"!��N��F4T�y�#Z)�1.�>(�.�oŅ�0���9�>�d��JK����5��95��q`���V�G:טD�t<kb����i�����~�g��a].�Ĉ�0�B�#�p�R�{OE�Y��T�=��ͩ��=!��H�%� 1�֞�0c'��+���؏f�V��x�'�m���]���@�\���z��z�ur�pc��X��E=	B1���i�z���nQi�2��P��H	�M;�+���JZ꯷��گGP��K�I��ș��OF�_�I�&(��6�+�4i:ox��������k�"�o{"�6Y��n<�m�T����>��N�rU��*7�,u����f����?O�vv	�;�vJD9���z���-�Ųk)�����Z�WBf���U�yOL��AS5+\��:����v�1�78v�`n��Wq���d����'	��bq4��F���b�DD��:�ݝJW�9!#�V�h�I^mر�3	gJ�4�ZDR[��{��#�!FX�%�*XxX����s��?�٪��Mp���`o���@:l⷗��(��.�P�h�>dc�0Z�3��Y�]
:��2�,�yx�ex�}�����Yl��/�{�Mȸ���q2���. %��ޑ �����[�ˮ�,�j�Y�p��{=.c�e�N���ꤑ��EQ�#�M�T��r�:�+=6����a5��z0�x?�Y�T�N]k]e�v��eA-��O��u��*:��}���j(JG43k�ލ�'���Ù2E��=���~�V�a8�L
֌��X6_��!�|���B|'�[H���r>�Dnv�Y��Yz�`InFDn���7�O�ר5�t��>�8��-{���#�HW)���?�� .�Q��ΜV��������c�:�j�s�����n=�3����y�o��Yґ�rO[�rVy*��bЕ��tB�w�i^MzA��l_=1!WE�8G�:J�?t;�'�X.I>�dj���� �G��܉��'P�3)���O\bs��;U�(�}x���1������n��f)���7i;�!d��:��j����f����唐���ԓƌ��^~c�� u1�r�6EU���2��Ƨ3�A��G��� 㩟��l������!}D��T�3�sq���ޡ"����Vu���V3KϑB��fŐ.������n�Aٴ�����?�����D�lS�Dv����w��X�JЁ�'��A��+uO��Z/�� ^�ݪG���:zX�E�8ѓ��Gs�96����<{@|%���As1y8��V�/�
�f��H[��}��"ƳC�4Pq覆�����z�>������<31��;��/3���j��HH�P��o�qe��ˎU�Jh��}���4_���e��m�.��J$#mv���7c>��5x�rh��:��@�v��QO�ؔh^��;<%���}2�8dTx��e�CiqY<����