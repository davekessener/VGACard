XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����b��và>�1���N>���6'aH��ked� �LN��ۯ,�}rA�}yS#����My.�y{�Iæ=�ڛJ�A�}y�L�]66��/�S������n�Sk��b���e��CQ��6�ޮ�W������r�*OH�=���a��_�9�k��ލc�Aκ�i�����M�C���P	�qa6�Z������B��T��5y��28�c4��$�Q� �&a��:x��D
��VU�c���c��n�Y o'���)�� I�Ͷ?17ù��M����2�8�>�������^ ۝�$X1�z�����JS��a_�1C=FR�y.�la��g��!����;�a�_� ���z�^���>7�]Ԍa�����l�����z,��Nw_��8/\(A�P�E���/�9L%2��R�}�����p"�!�cj}a�cGV�#����<L�����
v�do���[���p��g�i�k��=9`���δ^� �Z0,��-���2�k��!a�(��?�)�X�]�O���Ä\���=��i�+.�cjM����i��\��3>][́�P�h��F���Ӕ��>О<9����1��Y�[x����@w����&�7������q+ ��&e�	�4K4yݝ\��h�-��t�z����	k-g�OE@�ç����@"�o
�7�ޜz�-���1�4�$%y�/h��c�dQ��χ��Җ]�����k>�usX��c�y�����!)����6�{KX����XlxVHYEB    33bd     c90<��L^M���^�����V
��[��vJ���x��ٿ�Iqyy7���-8�&�$���;����&����'�l'5�l�g�!{	�U*)�,㡋H����U����F3Y$�c�rto�+16.�)���Bs�E�nX��#hU�c�������.��^��E^�S�TG�(�d�0��UN�"�/�.�-�x�y��韍\7�{&48_#`�lc#d����'�R�������ǂ]�d���o����㹎��	��������	�Z���+��
���cZ�8.��� ��1�酪T4��/u�{O �����������\s�Ө���!��	�v���*�� m�&M��ϏƂ�X�x`"�0�..�̖�<1��~�iS;1���fc�2 �?��#2#�f��L���^%�رRzm���l�3$�b�b�{Po59[R�@��ų��:��ӚX���Mh�`ڮQ��)k��)��a~��`:��-�*��9��nz��4�̋�QS�E���D\�����h��]n��E�8ݭ��h�F�C�'F.��o�)�@*j��[d��_N��	BrxB z\[�	V)�ލ�3�]MǤ�)��$�(`�±�WS�8�uA~ {���E������	_�<�����ѺVȰe[~�k����?�a�^�Z
~�Tn�x��Z�X��;󈳧J�DZ&�ZA뷴#��
ż3��M>/E��#��������*cH2��ä����>�a���t�]�3�,;_ql�7���w>c��yi�X;��+��-�I���:C鲋�����_P�U澚0����X=�zh�1��>kr#Բ��n䚚P�o˷�1��(�CBO`o�)���D*�e�tM�2�k!}���*
>t�\<�&
��&f�TmP�1���_s���%ih`�CI#x��Y��W�V3��fj^"�;@�y�я�b>�ԇ�<Y��{�� �|^��4���pck*FIev���vo<�־.9q E��A_H9����8���F���b���؜:{/r,	y��9�����}Y�����1ژ7V[9M�c�]�YJj�����p/JX֝�v�$#n'R� ݓa�#	�3�e��W���Ǝ�y�sĸ�sC��7�/ ��9�-�j����AYl`�60V���Z���N���#Ԥ��K·1S����4��=?�(Unpxb���N��YI��ޥ,̸��������X��D8�ݑ�d
��gNi\�p�t�HNb�'w�No��c ����{z>�^�{W�y�x@�[��3�	J��Q����R-A����@����We�kV��Ō�szE>��h��3!�^/F5�EE������'�*���/��a��I8��s��oA�s��C���f��ˑ��;��a�ѧd�v���6�x�pⓘʲ��9��������}TEB�l�u2���X� W�O�k��w���c��8���L��������pbWG�.J�J΁WzmRj�Ӳ�DS�c/�v��ٻ)��:�k�ʘed=�M/H��l޷�	�4����\圲�$�dr��N�O~�Ke��T-P�C�с9�y�N�����BL�*F��W(��x�N��[�C��ch�3���QHezvJ�Ӹ�WWռ��Ɠ&�vZ(=��Ëew�<�(��+�
��"g6�`v)C�� �n{ԉ1g�=���jա�a �,������Ěy���E0	�B
�F�KB$Rݬhi!�\�+���&`9�>��%΅��F+�/���� i�tz�"Y��ym���T�)7�'9��X���V I��C�>�TG<V��mynk���(�ʑܯj���h��:4g;�jd��K ��^K��d��My�`_-8�> ���m-�>A҆���	���7{:�	�0FN�k���03[x�8��k�*1����&#��������`ԅi�׼5��s��ֵ�L[+$jv��͑Ƥ�f���Q��3�5���@%Pu�������K˲_�Pȷ�ڈ�:͕���L;	�qv0��ˢ���m�n\x�A<+�R\k%�;��_��wrPhq�2�x���]�iG�V�-���(ަNq=��� �	�|	��6���r�6�N�RR��b'�i�[)�m���7��Ϧ������Ȣ7��J��/��.��)�Zk6�1�R� ���a\� 6�$��QF]RuwG�!���9���y��[�xL�?�Ԛ(m��p�cI^��hi.��R����-��ɋx����Y��J�\���	)��M���(�:���-��N���n��b��RY�]�B4�sWV	U�;$3�9W%���Jߝ��?�;q�q����U�j����'��n�gC�38(�%�s�)V���!u��_J'��x�	��:j}06��6đC!0����b)�͹�a: i)1@'�J���䇨�xJ�w�n_i�4�P�@|�@	���j���u�̴o�-Պ� �{J��u|�p�4M�{�J�����g2q�5:Rϔ���ȶ��g4i�/?jx#����w��'����j�r H	��"������I��:+>��-�h���������XW���~�8 �l���gm $�a��g�GdM,����q�H��+7�b���]J���T�*㚴�[�[��R���)[0Ph�l ���`���>�b,���q���m�&�5���%=�I�5z̟�j+c�K�qAvkP����[�D<���K	�?,��	 ��!f�y8�����+�8���gP_e�ƉS; �Ҽ	�pM������r�L�`>�iʜO �z��Yi�Є̟|��6�<������bZ��OM�$�8��x��P�q�Dc���qtp���xO	ǖ0d��	�n+c��̆3��1(Of�==�F�oX5��鄂��<���]j����ȃ&|����$�#�(����/F���)6���v�(&��1�!�_=�f�R��O��'�jE��i
�38�vj�{��Kϯ[m�Yu�ڰ�Z˅���ۤML�mB��c!/� �m>�
����M�	Zч�-���]V��EpEum��M���O!
w�bāB��؅r�6�s�qe�	�
�!OV��9�0���1a�v�5!�g���6�kEF��?D^2(�j��1��\���dZ�����U���9d�3�jH����e=�t�F