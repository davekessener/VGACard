XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���y\�$%�0��3�'�r^6<���S���oӌtS�Zs%:�ąyFގ����>�7�K1��&|$�w.��/q�0V?�_:v��p��%����ɨ����2�fU[��ɾR�'�S�����E�K��}z<W�[�UѸ�YY�'�[�s�`��_+���4���wZ��t��㻮?V�MzZg%�\����;q�V�⤉>'�Q8Nb9���C����΃�T�����#1M�./��#�ƛs���(��M4U@�4���@>��/R<�������.*/+C��u(ߟ~j����"$�����u�F��YM�[35E����n��[�	�v�y��~
fg�'�,`�x/D�*�_�|���G@c�˗��J���OB�Ȁ!�h��_,�[�$�	�5����q0��v�����/�:���f����|���,Z��-ڙFF��ᗹ�1_|{�Fl[8����Y $!��oqδ�n4���ܝK�#Ͽ�AO`���{~xp��ћ~@��Ӥ���p?փ|�CHrmX�W E��W/�I���BӋ��8�v�Ϗ�0퉞�o:���\��K2F�Xf:u^Ns���N������Pglͬ.6��'��q,�X� �I�.D� [���h��zf��'���P /q\�`i1�UI�ʾ�c�d���Y���a�mL��k�:������f-� ��q/JQ�
�>�3{l�e�Z��_ajG��3F�����
q�;@�㉐�/��W5��y�n�XlxVHYEB    b631    1a00bjW�E�� �ر������z��c�җJMj�[vbS?�>=a�9 ]Q�~���}�����'���?+L��5d�\rp�脰׊G�2�,��ogy��AeMX�z����'2G%�FZt �v�6�]�P�B�̡��3&LL���C{�	Z�(�$S��)�9ܿ��K�R�h��Q��i]&��d�^�}`�p���ӊ��o-!m�1�,ћ��&��L�8�f�M�*��&F���o�/^
���y��Q8�?w�:���EU5x���ޯD�I���*J�����Xh���P����8�A�E��cv�(j3>�q+R��q�����>�X>��$�Y	�]U��RFB��pyNޮEM	�V�}����&j���Q�K����`��!�6����1�hq4qb�#�|�<$��n��k{%�VP�.�T��X��Nx8�l?���5���m�y�G wȀ!��A-S���h \@`�+щ���[~{S��N����	ѹ�!�&g��$�H�]*K���y8W����Ԣ{��g��&g��t�-�1z)JHn�&�'up��b�Y��I��~K��������DKS�t]���*��DL�����	6����^���^~Y�ʘ�rA��x�_�U��GA�9M�����l��H�]�83����	�J�Wf��<���F/�Y�v�[�l ���V�Z��^4�֒���Ɠ(�u�Eڨzt��B~~��=8��Wh�~��D���k_m�L|<��ߍ-M��	y�ӈ�Jn�p+�w�l�t��[!<ܙ��r�7̒4����������~�-�a3��Z/F�-��=۸vA1�����/��@�L��T�'+�b��!pHsY2���31hj���͇Z���8m����1�D�iS�Q&�M��'[�������	(3��(<ψ��n���H�j��B�q�5Rɖ��/;����~�p�V?�(i�! :��*u.���AS�}>~5���Eif�+�]u�V�ɡ�N�����LA�:4���xa�ɋ{� �yI�bwH�B%���Qd�{t�����ټE<s����JJ�%��Ai\C��� +��OKGbE����[6'L�������~�}�m�IՈ�ע��	���v�a�n]��~�J�&��z;��i��O0���Fm�R����$�j��"/����r���nƏ� �m��Q���<�飔d���9`����}4w ��]=N���,F�	kein���X�8���SSE��j#^N�*�QM�y����v��ҟ~�rr�`���	.f�?U�x�\��{����bx�6�u�:�Ik��- "<ŷ-2�/d~kv]��� R{JU|{��l�����3>�jf~���ਫ	יW��Y�ϖ쑬.4T��r �E37$�Bf�Ʈ����e���=�%SWgr7���� }��c/Щ�],7�Wهx�uZ��/q��\0��S�,�mOQ��a���_�g�y�������^�t<]�A������[��Hɤ���)T}���=~.��v�<��"s?��&��@lp]lN�8����O����+�#᤮�%߭���f�".��k���5����p�N@�N��L��״.wr�.���]���IzP~��6c��@�4ɧ�S���Ԙ� U�����G�,i���{H����ߔ�%�n��K��!��a�`�-#4�1��Ժ|�q��"�,�︈�7ܚ\n ��1������V��h���JY��~ou��+D�	z$�I+Èl�'BX '(��Yh��-f{����9�g�2�B=�d?.l�I���Dޓ�o^�ƾ�3���#��&3!^�X��`:�C�zD-u所!@$�Z��]w��
�:����9�w5RS�[M�e�]���Qa�9�8B����V�����@��$�t���eI�|��Н�(�������Y��G���Z��b(wOHͩ�dp��J��t[�>%��ּz��N���-���=i��e�Bq��5�Ϩ[9i�a՚�Gw!���H�����ԃ��.`���/r����q4��[�R �����_aff�V�Q��pP&䳒8Y��`�7��_�`���	K.�R�6�"�!"���i#�l�E�n
B��q�[�滥���8���i�Ͱ)	I\���R>e]���3*��Sh����X�)D~���1$�b&E��P$=�Ώ�U2��Jm��g�5#Z��#ܩ��&��սxNA?����^�ҰCzZ��R�.�-� ��He������t[�_��"/L�s-C�k��R� P'�9����QFqL�y�L��g�D�U.-Jvl\�|�Ŝ��ԫ���&��C� ��P+&䠖��8���(,1%�k ��[����A~?�@ah��S���K��4�E�^!��o���Yy-���1m'���0��.,5�U�8G��k�m+�wծs,���O&|���$��%�o�ō�$�#��hi�8�E|�lQ������U��r%�����6|�}���/� z>�|�:�ņ�] ˼�6�t�"�҅ ���ө�C��1/���
K���WQ\�?��g��,�� �y��{��Ӫ�/���0�J]��wV_J�� ��!�kd�5��P�y�`�ijJA�R҉���k���wc��ϫ��1P�^����X54=����6��硠}���r���`�Jp�6.VbN�|6|��͓_Լ��)�x��	�a���s�Tw�=�tE�9_C�AB���S�?~�c�1�7���w�k@(6l��8��th2%��ʕ筍Fj��c9����%�7LP��+�c�Zv���-���?�_NɊC�at���kw	Ju��K2��ׯU�QJ�sb�}�}�_k��!�!&��8MnG���zqS�4��g>��y|0U��;���j�4rV��x�a�v�	��4��jbM���"<�|$E�b�k�����ZD:�<��Ҝ�J�H����n�K����eUɒ��A0"��������ǌ��}�W2�f"�Z�@��Y��:�z�k�|�=舑�����_�-�����u3&���e����8�=��	 e=KNVj3Q��:�=S`�|iA��;�k�k��r�D����=�9��������*Ej}��3����R�]������DGN=�[7��/�$,��?��#��2J8'r�S~�к&���k����#A��$��O�c�?�:*=6رvr�%�$^�F��K�ޚ�{�����X�{����}��g<Ž�;B��%���V�]F�#b3:T�|�e�5�Έ�[��@��+ٝ�5Kf<" �t	4����W�!w�g���Uw<� �(��)���yC?/I
�T���e��N�_\"��BJb����вG�pP�7��� d *�"��#�"���v�a���*3���o��d��F�	%�:�5���~ �9��a8���ОBe/SJѦ��c�+�=�Ӣ��/�{�b�[f����b�8�c�6��mK:h�JeTDU��h)-u����7�G�@�q��A��Mir�EuhPr���b6>,Q���/�ӑ$h�!���a`�&2�DH�>�I��?�1�-|x�iU�A��2��C] �����g���f^��dX�Y�Ȍ����f� �G��wf��c���ɇ�6v���^�e&��Z����O��'��GUs��VI�g�`����:��.���Q��ͩ��Nc%���L,����Ў�֊���'�b�ʆ����M��^ޡW$��X��DJ��x�Y�f�P�SKhc+����6XF�Z�s�C>��P�7����o`�O�6�j�����t`�m 8Z�zK�^nu�f�:Ei�_�kY��U��.8�h�Ѩ���8��W���dC�x�i.��K��>c�;,�-v�E{�1�%�I�g��'�`������!�g�u������0G��6`2g���%�@�O+��]����e��^A��P���d�in�7Z�
��H 4�w*.)$���#+��qL{?}NҞ����.[�r�
����6�O����y�Ї����H�W�
���h�Q��X�4��D;.��^�z�2�@��X<�g�3��ѝ#֑��_1*��������}��@q�;�����*���w�uV��\D�O ��3�HoE��!��dޖ�*9Ɍ���>yDR&h� �abV��3�R��Vb%4@ci��x:�����aoʖ|D�Kf�yϔ����,���s�S�}��Ae���,x΢`ݻs����ʑ��6�	Y�2��(��K�AO�ץ�ƅ�����a�>vfO�Z�Y�%��}AHVu:E�u�	?� ��N>�c���Mg�DK������_ES$Om|_Ő�~���Ծf�$����D��j�
����� U�.���4~k:=�k	���e�ԉy\o~)b�H��Gx����Ye�<�o�)nf����4��k΅�A���D���ҋ��/80clVz7b��?�)��W3E]�78-�[s����5�lY}�,��F����y��n[`z��v��a��c쾱x�5�%�t�M��jZ�������!�u_��&�[n�Y�����å��cr��n���8i�++�r�'���N9"UE��9���R�;ۈ�&m��
�R��Ԋ�$�L�Mӱ���-T��+�3=�"�<W������y���~�7��0o�y�!,���>v߉��` f�z�����l��BM��9�z��Ch�����H���{N�I�#���sġ�/�]�eaMaI�$�>62��Qn?�{�'}F�3$��l>�h�X�dy�F�m���Lx�W�@R�tv8O�O
�����6\�p�c�q���󂻱�
��,ד������G��͛B$��ELږt�Ry�Qk�v�$�`���dP����n�e-�0<�v�lg�g���8��$<8=N��;; �K��Ԩ���Q���s�җSeN��͠l��j'�k����!!g�_]4���Ȝ��rt�
�CB�d����kg��G��^~𗶏H������p!��NqL��;�����%�]�?�4��}�Tl���!7��0�8ϙ�����(D��mڴ�u�Ywg���-9���lp0H���H'�E�BR��_��M���*N���:��"�{p�b�G��k��������<4K�=֍\�{)�Uqh
'����Mq 
���op˟>�hH���A�vI!���\�xV���	%� >�-���}�[�ml_�i-9�*e&��ȇ�.�'��	+GR���;�cq}����r�d+ R�4�Ѫԁq�>�9�Xn�or����Y���`a4��Ͻ;�x�?P��E��O,V6� Ch���Ō�K�����aU���B^x�Z.��zG�zT5f�t	]�v_ϯ5�B=���xjr����>7�J�y-��fW����@�ڮ��)�=���{��Kh�9�^�K�E����7�s�v��lrN���/�������-���?��rtڍ��i���d�� ;ʿGzr��_D!Ǽ]W5�J`oc�:�Eaaq,8c��Uh:����@�~\����u�+�D�4�������|^*����g�'s=����wL���޸=B��ϩ,ե�"VFt���)�#\3���=�Xs�Iߪc�w��;%���
f���[�|��);�omR�{^�ݣ���f7���7D~�ٹN�V%�]�$ٖ���%Px!Lš�pp@JQ�>�g�ٷ�JE�FA��ʹ��ȣ�g�/|p�SR;����L;�@��)c�kqE	D�N���K����W�<�<��>U%˻lB����������W�y��������L��f����I ���CHZY �d}"���'�\�odg�\x&8��\kY���۽��b�tĔ`Ϳĥ��mVEE8����K�"#���X�Γh��J7A?���+����g �[���g�xr�H���Ⱦ�T�}k��?��&n8���tV��n�c7�F���(en�+OM}ѵ��\�"�U$
�RH�p��q�������2@�XN�_�s/T�{�b?Z^z�b�����l�L���͌�-������4:�r=PGOWS��b%�V�@8(�{��
�o+��{�Cf��*m�A�&H���	� ��4�l�E�cR[F_g.K���淔����|��5����h9��z���	2̛�z6��a�v_9L�|)q۫Hn{b��`��Đ�
���/��r6��v��W�'%�>�PZi
��Xl]��C� ߐ�4$N��Xa�:�I��֫,Q�_�Z i٣TѬ/�d��t��mB�̪��Y�%���
���WH�v�T�ۍ��ĀU.|��^�)ah�zK~ީGD��V0#����*��yƉ<���:?6z����Q�E9:z���78�Y�	/���6۹���Z�,�@���&}{di��z���n�X�X��[2lg<_������s?C$J��<�`gfS�͉KuN���]�Z��A�xl6�(�y���Y�-��U�!���4������|p