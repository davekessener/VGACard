XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���D���y������uuσa�ɱ(���ȝvS..�2M�����=�������I����1�4�XȰh'zv7�c)��KOr.�hȇ��z��HE��t�ʇ��_�AIM	;�D�yZR�u��f�� �Ӿ����cD*�b�"sBb����ۯ�$��(���j�ܧ��3#��Q�%��-^��<~�g�fj�qw����UES<N�����//�f�g�����բ�pq鰅a�z�2Q�_,�Y�����qjY1D`t����B��|VV<��'	h��tEs�a&ػ������q�<JC�Xb�u�m�_��vK�ZCN)2s���+E*T`tS�ۅ��PF=iT
��M1�L~V���y^�1����̥حG�l�[�dO? �L
��lr�Q_�&yN	�#�M4<�U��ӃZ�D�sa�V�h|{��Sd�;c���Z��w(�Qɚ7����	&�T7.0���}	����˞�[f~�pr�c��~�i)+VH�M����7�DDw�x9/?IT�M��b��OZ��ky��n�7�-�T���#�J$�>s�w/_	�(qVWVT}4��b�Bg0/Q�%�� �?��kA���mx�-�֦H\V�� E�+��'�G����A��Z���"N1^Z��|�����D1(�u ��lb��a�n�#�hи�M&ؾn�7g�P��>{I���G���0B��L�e:�ڝĔS�����su#�`TMr����^�&<���P�����#("�I.XlxVHYEB    fa00    1950
��hb�@Nx�s�{b�A���(!�̛t�I
�U�Yն�+�Ϩ3+��O��ײ��Abv���H���U��3w��i��q��%:>�%�׽���s+<��W��0�X0k��ؔ�h��Ĵ"V�j��f��K���>����G�B�����q0T��d��	\i�ʌ�A֌o��!(�2z4��n*��G�坁��qc.،�ڒRH`i�{�U���;�뜪I��1B�n=�?��Ӱ|05�ѪG�U`�fdhlif0!z���V�Q}�ᔡ�y��x�XtQ�=t�1'�N o���-u�P�%Է�΋��l|4�ѯ��b4.�����+�u~W�c�;w����Ǒ̖�Fi��=�b͚�t%s�ׯ�m����<mI�j�����Zj�::��}�.��m�S�,V}�R[��-�#PN�r��f�����`0��C?Ciw��=F/q'8k�q[�Y�F��	�Q[ǯ����i=��ώaO���-S�ȉ��b�+g�R������'�RȽ$t6�.nqm�w4�.M��t���wdx�:�j`���#nb��EKŌ<4�Jtٕȡ��,kv��ڍr��F#Ɯ{tjR� ň��M��xD�&�M���}L�+p�ǧ��,,x�H8a�[ ��ȸ��\��Y��#�o���.��*�f�(���5�xG��0$KUMK#ٿ6dT���wR�!
�&	�jFS��Fȳ��$�s�5�i�L��ˉD�\����**�ə��ϗ�)@9W��g_]d�ᡄ����-���g ��o���D�H�9��cek�8���Y�=�3��e	�pk���@B�y�d�<b��w&UtL��D��q�W�S$'5�6q�pυ�W�ea�^��.����g�����^7���٥��sB2��]�n�%c�1!6cͯK��Q6�p#yq�E���	�NR8ɞ�ƶĹ���R�q<v&����s������^ԄRi����D�*B���BP���(|&�D��[��rE�r_|��eL��n����iA���M�=Z@��ɟE�^us�5�D����~,�F��+M��J��
��MWV��E�+�	J�B�3Q�C�<U�(O�s�c�\3y�O*�N�d��z�|��}��$��9���w�v�zG�����pz�	Y��`�W:�RS������P���y�K��t1���Zx�5���	�<���oEC��/�K����I���Ʊ�^���X��\p�d��CZqHe���[�$m�5��U��RJq���xUh�|.��F���=l�[�I�%���B[��S7�#�_X���Vgm��+~��jL &X�h���M@0���W6$.��~z�Dے�ar"��뿨�F�9�z�(�Pͼ�پ"��5�o��S���s�����{]��(�B|Ɲ���1��!]7I��-ŤjF2�M"Lq��n�;?��z�l�P��)'$2n�$�ۆ� ��V��i����6�j�����<�������J�g���o1>*_&����KK�p{���/j�& @V2�P-�l���I��z�<Z�L�[e�.�S�����.`ddߊ�n7���`�ce{b�(c!1<��������u�@�L��9"9�=\��gHUB�������Bo?p��o�4�*bv2xi�g DB��|>���_,�fL�m`�D��c-�zsp��r ����m4a�zW�j���o�;�������FSJ���"�d,�Z��O�>�b�I9p�(
��M��)�W����!�:{^uR�3c���~Y��Z*L����(G�FMr��h�g�bnbJ"���yvu�,m���Yǲ�c��р���Rζ� ��8�~��P��OD�%�
�b�ck#��^\p.��D1�oZ6XY_�l�����[Q��ZFPy�����ړk[2�]�)���mD��XW��2�m%+��[�Y�� wzS��\sĒj������~2G"�,QN�*S���%9@����8C�*�ؽ�3��(�58�4�p�������Nq@�����	���>}�K���3��v����3��X�-_�0���R��o�|��Q�u�!��ң�l!��F$K�ԃGG+eg��ĈH�� ��qi	�I�ӭ&A�C���;c
\���@����B��J��!�Z�6��Ӹ��sLR�:W�oc�=��v�@8�K���Q��+p��ԥ�*�l��vn�^n	GCE�,�R6��[�`�Oe�FP�p(&忿p0�����c����iQڿ�U��d@�؅��;�8R��sWm���n��6�{�/vA�;w��<����L�=�t޼�� �ufZ��E�����(��nb�u#e�~|cq|��hVs�Bdqj�!5���Q�h/Z�����Ha��Ʀ����2��?��}b02v(���9�rXr�^�&��xz�P_�ӆ9e�1LX�H��Ho��>�P�^g+��tLֿ�p�r���"��W�B'�=��y�n���D�Z��hrk�Y�wl��~���:�a��hǟ�o�Ե�%��_p�*�n�'��[������h���Ε�8h�iL�d�7y�<N���
��&4����*�P)��A��P�:f��L�Gp���i\�`rEs���I������z��}vsͱ�9���?�!�`��\��}�L�t�sN��$&�����|��	9]���1>�i/���9CxN����/��(4�F���ƥkB!#��d/����+xs	���h��. Ƨu6p��:�
>̅]�lQZ0����	`]M����/�]�P�^NO���ui����¡G�iһp�:鰘����`�螻A�h�!�ۻ��p�/���OX]�嚃���X���]]m5c�j ������N�g(P��6#�X�ŵ�d��u}�XSԩ����ݴ� �*ը#2�ԥq�~MU�����%y�ŝ��"��}7����Y(�Vĺ��&�RX8'��Ů�oͷ+�@ksQO2s����<�������o��@+ܹF�qs1+_����6G��O�Ӑ^f��4�<ۗq]�w�����0hV��AM�y%39�
�xk���zѷT��:�n�2�+����oK�VB��p��f��11����2����RW~�L)�]��O\��:f,�]����$V���l��k&3�3۠���`%�/"1��t��s����Ql�u��jW�@�h',����2�|l �PqD�Z�K�H6��%��c!�9�xjYj-i�Zϴ3�7�������j�z H�>���	�:�T-����}���̺F�|�9�SRV�J��.өJ��կp�n��j�͒n��b�uķF��5!�\'�w�ݪ5h���n���-5:9DV��C�[}�[�����ì��"���ws��I��,%ki�
���b��g��\<�fz?��^g��ښ�����z��PF!�����5���5�uui�q.ߩM����Io������k�ᴡG���J����˩�@��pd[����n��m�������{I�´)O-0�]%����Լ����4V���ri!v�0��$R���nL�%p�6V�*۫A�������� ֳ7��N���,��ڟ�T��B�:~%,x�@+��φfG��r"����լ���@D-��j.m�\� ʈj�VƼ�}�T%ߕ6H%��,��+�92��gD��w�B�`�u�k���^��z�.k|-=����i7���T���$Y�J_g&��
��u���Y˶g	��-����33���Ƌ���!]�}��/�<�#tU}�m�k�P)�f$8�����O��T��]T0603���Sg��3P
�^���=����9md���Z~E���{6�/ıF� �E�˟����C�ё�J;���[�;u��� ��4S8l͡�J�G:8G'/F��T��)V����:tɜEqy�X���A�5	��)�r��d ��!�v���=΅��s�n^�#����ge��2c�1m��հj���i�N�E������ �8����%ܩ�\/$ZI4\�nC&`�f��^5��"s�.ܧ���AD��y~Y�8�ڙq���AR|�0�1�Q=���e(s<��MIU�XXB�-�K��!}3�3����)�N p�|w&�fzI��[(Us`w��S��-��dw�5�b�7
��V .���>��O知��3��\�K�YS�?�̞���Ae����66��0Hr|�̵����Bp�ޗ�2�ʁ���.�5���M�`Ks�y�>(Q���i_0��/7
(����'x^�)� m�)�k�cz�����Ue�;��u�#��cI�~y,���b�uR�So�P�,�����
+�:bC?7� G�z��g�Ϡ�v��b�%iYa�o�:}s�1����s{��Ǘ���mr��"X���܃���7�ka;k�d)�|X��uȠj��9���j���SpGc}N�Ӌ�������IE��G�<�]!Å�OV~���cjnU`;���@2���`ԕ�J�RB�@u�ϣ$������E|i�B�k]��&�!�|c��r~;T��k8 ��LǏ��E�p�O}�\$j+ Kj�qKl���[�&�Ze����	v�.�Ŏ=�FD�u_�J�e�� �pQ�E��#�E�ꅨ�YF���p�MO5��EVg46x8�M�!���vh����aH�(ۨ�if��I'U�t(��5Sټ�c/n� T���T�����۾��)}C)�t-�PCY�u��G�3Ǯ3���x�����dB5+hkZ�����ԟ	2ȏ{[�J�YC_�ۋK����n9�x���l���%8p�;$r-a
���vSP�A	�
��?����&T|�	���G�%�6����}r���GuB�l���uR�TI��g�`�C�8�%��ɤ�U���lk���vY M�+�y�A�ֈ�?���m���1���ZUN��2c��s��y٭�PŴY}���{���E�����үs<Q�^���5oT�����T<.���f��e��mU���)�,@��5�Ue��/�7�o�%3^|i\����.�\Ȓإ�4�l�"�BCX"�%�������ЉN�Nx�Gz�������-���5$�0�����?�Pq�'��M�dB��)k6�[�fj�R2��2���	����!�!rft8=n�h o�u��g�rLK�SDvQ:�p��*c������m��G*��k�}�ӗ�|���ފp�'�o6�|z�E�) 0:@��;Ͱ���d�{��/�|pƜٞ:��d7�CY\���H��qۢ%���Wj�vk@s���0��,5�R�؛�T�^Җ������D!�F� Qn�?��G�n\�"��#�M�o�-�nz_QNgIN���~'i��� ��[���'�F�L�Ǫۡ/��"C�&i���1]P��U%)l�cU'5H�,+7��J�Z��4�C�M�
Z��{���j�'����7���,7'Jx�VJ�離B�o���\"<l�2�Y�,���'~+u�9�ZW���+BzL�Օ�T��l�5����L}�(ʗgv?C��&uh��Y�~�O]��>��ku|�6�1GK��V�ZFj�vu]��$+��h$[�
{J	5-�E�!fؾ �y���*Td��_(���f�.x?�(�%S�%@��zρ�g9�^v)LO4�D�w�G�y�N����M	�k����g��̆=G.�1$YN�F���X^�Bt�y��}c��ɀ�]f�T0���+��ٖu8�����74��a�`�  �_z����=OIR�a�W!Fy���(�A6���ogk����6=�?U�$��ӌy�E3 ���R	ƣy5���g�h;��ɷF�b��hҰ���'�ך�XyO���%ǔ`-T��]�
bS�o���͋DE|��ЅK�Ӷ�m������,e$R�;	�,�R�dPl����q�����S ~\Y�~�w�f���Ύ��:-��D<r����/��}��H� S��M8��mni�����v���.����k�Cs^n&:E-u��k�E7�mg�1h�ol��t�+$��{���5��?wXd�#�r��=s�D�'�Ƈ�n9��vF�F�,�h8�����b3Dv��^fV>�.��5��*Ж:���?V#�]V�6�#�E[��(��M��&3�悏�WVw������S� :X�V��Xv�!-<z������zt�9��%bj;1mQO�~5s�h@��c����o�ā��2Z�m4u����qH?2	[����)H=���'��C���W�R�Yw�X_1�l�����9-< c^��TNЄ[�%�3x���d5���|��Or�gKfnV�\<�� c��x�9�p8{����UQf����Qřۋ� ��K��m�쵇KFzҌ���u��F�ԔcȒ+P�XlxVHYEB    fa00     700H�c���W¶�wj4�;_'�P��wC?�X�5�"3��'b�x_���U`t�Q�:l˵Kv�1��~�����vV.Y$�J��N^\^�fEQ@�%,G�*��W[���y��{�KE]�c������#h�ȵ���W���kL�.��0�}}\_5�/^��D��I���HK�&��etǐ�~�:�L WR{'�A�w~����5M8%�M��.��흉�]����C/�m���荙�5�v6��(�C�%n�݊[?]� ��V
��MF_�T)��j�EvbDG��*�e��.Yh�����
Uv�(��7�eg$���K�ȳ����MJ\>=M 
��9�x'���U�kq�,���SB)Ӎ��~'Ƭ����4��#��T��b��%z>n��(��W�<-S-�O#i�s�T�,�:TC��&:'��?� z�˴���W�nq^��ng&����<�[0o�y�+a�s�-׺���G>�\�r�P�wD:�Xx��0R����Up c��rC ���~�cu'"BƆ��Y�j9���S4��jg�gT��na��R:%*�{��`z��O�����S9b�E��qR/Xx@_ˉ-�6��&0D���`���"�ə=��"4�H�0A���9w|,I���?�/ז;=/�	s�Z�����8]6͚2Qxrπ�7���Uv ��: Q1b�M����LL�R�JEB�ӗqM�z�{�n��eF�ϳ�����ndg������Q���nJ�H��.c���a9P�w��T<���RjW�oRA.ң7�}	�Y��t�T���b�.��=�a��N�{��}�0�ļ�2�Ϊ��HV�t�1W�0�1 a�&�@���1�0)��P�l��D�Űœ6�JU��_���r����W�C���7C�µ�c��J9Ң2^NXO��E�_����4/%�=�x�}�`�D_����NϏkyV[�ű�s����Wd���/7{������Q-j!޹)=>?MfGt%!>m��u~]���k�^�T�q�W�Sa�rX�>wo����~�a �a�0V4?�;a�N�'���ƺ����7Q�G����&�
��9��j�@Y�KA��\e����z�;��L�5x/�W�߼^8^<��
���ȸ������w��N�n_�ۇ��������N{W��!�&��u"��zJtQu� �\��1�mv�//�^IlrR�%�@��K��%����Q�1�G�w�#f�'	�����چC;}n93s|(H�]9/3�n
#��/�
����"�Ǘ�R�yNB��2ol9+X^~d�r���q]l�����y�ۿ��]����K��c���Z��WK>n�;� �Ia=�޿|י��������H����4Y��ܹ�x�*���/5'���x��*���%Zo�a��&(�����a����Z򧊔Z�W/Z- k�XZ�<��xS���3����Y=��i�N|���A�M�qY�Kc�u`��k0�j]��{�O��Q���豢|C���R�=���Ӱ}.}gU5.h?N�	��7�������д���6 ��Xq��{^2a�9��� ��D���5�z�g���z�¦^�߄c�����4 '���P	d˫IXlw��wJ�a<mjoE�!j��<�Qr����^+?l���,���먈(!lXN1�CGDz���}�<e����N���@�|�(R!Դ鯝J��x���uXtD��xdpq$�8蘬>5�x�^T�����.j/&�F���Afp��)��m���]|�XlxVHYEB    77da     a60�j�/�CyH/�hUW5�β��\�2�yx�Q ��U8�]��J,\��p  ��k��H�GL��X����{�p�h��Yeiq���OKv�b�s�p�\�����& �����ߐ5T"t���R
3�~W
ij���F�����M�k	K �^b��>�y1����90�>L��_$�n
O>�T����Sdv����)�S<]�îl������ /���-���T`0��-���~T���� gqy�Z��b8�b�-*7�FJ�.n[�a��h?$1��"�i�=;i�wk�Z�����&�=�K��D/~߸�R�X��1��ޝ���}m�BfNx0�>�_s�T�3rS�:mo=���9v�m���7��k2�
�
�'�U	��$�\@����S���1��K�=��&��LrR�N�.�r��1b�5�	�Ϭ}����$�Md.�n��c-�^_�"�u|ݼ]������\���S�/�$bo�kM�#0+o��>"w����8;
ja�zĘ=�b����ۈ�7��kyo���<�Ɩ/���8i���ʜ�u[��D��[X~D�Rb+����cVݾ��z�2�^0e/�A�.xCe(�<���������w��|�u���~�����KXr'@-�������ND�ιٙQ$ʄA��[ޱ���0�O�{꠿s����]6"�<6��������������36j.������̡5�~�B��8����K�!6s�&��Ⱥ���{��U�4�R�r�*�e��E:���*��^��s�W�57x��UR�\�A��8�I�����I��X���L��Xp�\���>�ô�3��a�ţ���f������{����/���Pxsk��(�;�w�9Y�$�����7����M�~�mETσ��U! ̊d?�V|�O����I8��1�Q0f� 5y>�GV%3}ĭ��\U����Lc5����ڒxTсL����S�W���`�
��q�/�+��Y�`%7�d�=Ӭ����)DK�80n��� ?TOϕ����\1|�,Uハt	�xr�ȕ^՚�����-`��@E�����z)�`ϟ�eD�+#;H����;����#�"Е0��L��?����^iw��.� ���$m���\�d�v-)	u�����=U�Ώ�zj��hÑ��^Z�[n4Gd:�6/�:�
'.�4��*v��C�U&�_o�P81�X��ƺ�D�t�N���P�0ԫ���Y�/KY��v�.�G�����a��s�R�H�9��f<B�u��\�Ǜ:Х2����-s�2��,v��/�\X-C�\�9�;���N㑮"��r�{٧�鷃����D
`��R���G!����V�ZZ�nZ�r��K"���Ƶ��	��h��7@�^��b��Xc��/J�2BV��>�q��ՠ�����[i�Ω
n��k-��w�e����Ox�2X�!�fUIȳ�=�q��a�����3`J���L<m'�97c��-�)��'FN�Q�`�grխ�{-a���X��{Z�E�>$F�^�mLD������q8A1���sS�C�OSC�o��Cb�P�����'�~�[��J��D�S��\a`B~�~�d+�"�n��,�m.<�b�1��򧸈�Ppv�h�����5���Q���mpT���4n�5�ȱJe�{�1��ȼ��>�g�uE4"u���)����� 1\�g�ӊ/C�㐴B�(�>��a��R�%�����bc�e�1K�����o�ˢ��T�[� ,��,B��r3b��H�D�`�\ml�YZ�ڃ��L��ϰ�|�&軨kzb9�F�@q�� H����3C��r�д��ݟ*�f�9I'��[=�&Ku7���#��;}r+v����+�XU���a�~}���Mbט�0�q���VZ��� �Q7,�,h+gU�9u��p�jU?���^���|\KG/]�t}������)~g��&ҢjVɮ)��ɜ���Iڨ��c�vU";�c��u�e�j�b����c�}��o	�6��(��d��o%��&g�?�	)��8�d����#rľ/~xmI�Dރ��EFe�~ � �]�Z��	�Ơ�ʙQ�о�eެ:z���G8�"������f�"�ѕA��v�[n�Jܣ@]^`{��68��X�/�=��<�GP�(�?p{�^�оj�AĊ���� Wm�#���l��d9��J@*�d���?t7ʿ�fla��������XZ��o��V;>��r�If��Xtb��t]����.�5�Su�g��(����*z�4n���'���!h]�-��j&� ͜Qj{H�195	$��k	��xgVþ��u���yWs�]��l0}w�i낯�>��R�v��ځ�VK�e52��b���l�Cp��Wh+�q��-9Đ����E��1J0��h0Aܿ�i���ǋ�A�#�0��O+� ���y���,]?-\��L4�#FO)�瓦 �z�y/�S�� c����2H;E4�u8J�^ SƄ��f�>�=��V�V[p�� Ji��j��c�!���g(4<��>̜Z�ە�5��ϐ&��zy!����<��O+�a�~`oz��`���ֻ�,�	�Ϩߔ�Fõ�����!Z�7i��3�ű(JP��