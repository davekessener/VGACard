XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"v:���Z:��a.�i+(�tM�{Cɱ2����U-�#�!u
<G�w�hƟ2��x3�=fS�1}	��B��L�)���S�N��-7jU��޼_� �C�����|Hr��~{M�' X�,N���GX~2�Ɨ��uR��t<��<s2��]�A���ǒ��.��G7�-�0�C!��_[u�<ϡ$m�m?Q�D�7|=��y�x�WP]������-�;
KQ�,��d,�#���iIҺ[��r�av���]Nx`�b˦�G�H�V~O�Oa;�ԧ�.J+h�p2��%��#_������D<!��l�:Va&@�^j�/���A�~�h���{�"B�b1�5Gվ�3�3�=��Uz��ߚ��
Q��19g��\��1�ah'��� �|��}��{�1�5���'�蔂kd �Џ�cG������SBMG:����u���g��q������$B���1=��j�I��3i�{�\u��8b��f���j��ؗ�2���-l�f�W��K�1�֩|��#��v�ē}u2eJE;���$��s�t�,��K��QVZ*:a�2-��Z��D���B����RcH����j����i7�q���\� T���V_Z�>P�Ѯ�8Y��Q�}t�nr&�/�Z/��a����m8��4��Թ�Xִj������l_�
�8Bxܲ�N��Mj�<E91���7A��f0� �6SC��Q�J6Sg���,�B꒬�F��8��h
x�z�`T�Ow/]3�� �u-��Tk]_XlxVHYEB    fa00    2910s�9^�c˸%�F�ݨ�h�03���v���4��� ��lbq3�Q��t7�o��PqD�ϡ;�����
�)e�*��g� Oɰ����h?��	�98U3p�&�I6$�?c��A-���0�6K���6Mxb��,��&��	���+��[�sJ�*����n-��#�9?���YH��9$+ �m��RMN�T���V�>F�0h��>�O>��W�2��_�:IV�N����y燥r�����<��,j�<����h�į���z��y/}[A��}5>����&E�i��dR�t!�Yu)��Γ���3<���o��@?!���9�Ӵ����2�MQ�|HĄ�Շ���l�rQ���������U�z�|۲>�?��W���Q�> +�J��ͻ���b��J�/�b@��>��МqQr:\��t(�FM^�:�A�	���1J�0�A��tq���s�f�U���yŲ����5u@��"�qv�lk[���9'$����9�J��{�C�4k�G�*|d(�W*݊�,=�,�Je�RI��w�V���΃Z��a���K+�\�@�{�t[|����KC�P�8���x ��$f�	�^����cpxF89&V�	`�Z�㫯*�^dȶ�t"��{'�Rk꼀� P��|�R���UgX��c���]	�N�HQ�4��+�����W�bٖ�����%N��*�7�R3r=��. ��VB"�0��
��p0�=��E�m;�#a��Qe��3����x�g4��-^f��J�|i��YL��X:[<�m�́Ҁ]���h&Ba��V�K��|�l�Ġ��HHf+`Ta�o�%��EyU��e�oh�_�7u/q �]Mq�{�J�j���w��du�K#W�u`z�a."<l�Nd8	>��O��ѱ�3��V��Wk�I�Q
��q���|����3�K�}���u{���� �꠵�99�l^A�!{z[�B�$x�5��,��37�b��o���(�!�߷6����l<�gp�>�)ㄦ\�"ND@�7���v�7�� ������[�^jygnJ~��_�]����Z�w��j@4m�5aj�FN�9�
!�92�)�e��Ϝ 3a��	����X���K&��G'<-���G�Ec678�(nEL[-3����q�O?�����aT#����w\��B�\dC�5���if�L�}-��h�,��d�]p@ř`J͵w;���C�kpJ�`��I�0��o�xZ�rrK��4 ؍_��	FA�SS�=Z����Z�P�)��-pew�+�θ���ja�X2�d%C� `�L��<v�V���E�_��O}�(�g�<��k^�!\�GD���㆗L$����-}��o/0�c���|�?aX;��r# ��γñ��9�/�u]Cj1�D�vs����iEX���GZ�<D��kﵝpbJ#� ����Yj������O|U���/�`�>�����o�*5��L��MKf��c[�@�bX�mlA�#z���n��B���]�6wp�5���&5?CMVa��qU��(�q�,�2K��SE����S�^��4��Z�M�iO��U@���|�7�	��*3����U�W��AM��qT�:��񛱛,�nwF�H6LR�Μ�(�>�/2h3d�L��=�[�j�pmAsU�-��x���rh���(beg���U`�(�au�un���0��Ѱ�@F�1!>Y����ݫ��x��8�H�Ԭ%P�*k۠�D�H���ڊ�S	r�7�ͻ�!�pH�K|2�K=���2��M�:I����M!#{z�1�J�������(>M/Q7����ֺ
z�-�.p$��H6�zAE����^u����
��$f�]�IH�g���.N�Ϯ�F;���Z����4�i�R� ��/�Ȱ��T�W�2u���]c6�\�ʯO���Ca��@�Fp�]��|��#���P0�6[�(��J���͵4/�,t=�pw1~bٯ���|<C���o�dA�\�=��t�q�(㡦�ԁ�'3>�:��L�W���x�S��5���:xG�t�
,E�n8h�T3�?ʁ�=~2~�e��t�R4f�7�$�n,\��%��)b��q�<�����|�9���d�����
�
����$��j�ږa��סU��$hN�-Ԗ�l����xU11����Ѩl���S� g���*�aL�j�,^Z��&��-j�w
hNpy"���۷yY2H��J�@y��D$y�@��9�%��N��>�\/�ox�:�q����:�ϵm�A���fG����h�j؄�ͅ[�\i%N3w�x���i!A��N�8:xF�*�(/���qCй��b-sd�{5�%	W�0E�A�Jk��Ap�``>���?���଼ �q)��X0�x'��V
[|@�u]���#b�;D�xzP�@����#l�FLhQV}NK#�S����>d�dT��Ԙ����x�Wn-|�/�o��'�o��=d�=xl�z�2v����%���-��fA.�����n��91�3����[,�4Q�|����Wo��O�����r2L%A"�͌�=ZGZU(ߦ�x�?m�����t���"g_��i ��M�6�=��~)����X[0G�%�I'�����×��ʏ�3a�|EW�����R�:�DJ���_���랮P	\LufH��z�@��LM����nq�9��r��g}SЬw��I[�h�z���]�9���2&��Q��u���2x�G���E�IA+�<�1�DW~v����Ug+����(�4Q��X,�_�V���/�6�,9�8-�#��S�I��h�.�^����Wr�_�ן���^�P��Ri�y"a���z*c<׀�(9�é�VS�W��n(􀡯N�~���L��lh�/1�0=6?၌��ԦN����}V�D�"q��p�nH���-�j��'��>�D�=�'��P�KR��.��}C"�[ju�g���sۋR�ǵ��VG�T!�8s�e�-}=w}b֐f��$��cZ�AuC�T?����T��1x�p�6oy��ϫ��4)�"�j�4�l�;(\x�--�j�@Wv�h@�����bW�U�Ф������Hŵ#�_B��Sd�@B�9�|LzkM[.�x��	���g� �^X�3�6V�h��P	@�2�o7Jk~C	������}�u9"�:�F(o�����b�|�\���g~�7�f��
�����m�+�Q!�<�p�����aH�b�T���$�6v�;�~�!������8�j�|+[���&@��4/z-o%�|[��SL?/�	�B\��c"ܭ�xB=���l�D�-i���e�V�Ky�x��>��}T���៲�;�0}����8N�� u�oָ�C4��C�~�d�s��UyсՖ\�+Ӻ%В�2q���ѣ^���;񸯲C��p2��M�����~�1�ΊF)�jlب6�>��N�����[ؾ��������P7�o<o���B�h��h[��ə9�/M���^��?_��zӯ�R>��>���UAv��_o�H���^x�m� �R�g
~1��%�Hc73�,4_��ރ~�z�6�����$�}�5L�$�8M~�S��� �R�����g}���԰a�B�$������uY�12�˶N!v(d�u�)�I����w:=7{XӰ�f W�
3F=c��q�z7v($� �Ҟx��Y$!���uy~����\�Vc�o����]��Rz��_?MGo�-�ԓ�M�Qe^c��$!��vm1>Q�\�>�Q���̨��y:����ms��&6�0#㪵4WWj�#'����|a��p�g^�Y�j�9O�:��RT:�6�r�}-���Jm�DMDgN<�]N����ze]X��e6!�~*0��W�	��e��	}�iƜ���u�}|�F1 �M�M&�e�#:=��#!k`.�`��t77�s����G|��I[ZQ�L��-HWD�7Ӂ&~Hc�D���N�����7<3!<���̑$�ꚤ�P/���`���8hH�mIT�;��bΐ[�b'�]|F��c�i��n�;od?,V;����	��_� ��ǟ�.B[�}�����l3�"���
1�<1hM�q{��͛s���L-D�a�6�h���:�vj-�hHɡ�����2�_�~[K4+W�r�;H���:�P��ф��q ={�#:�jс2���D[��)��z�j:���`�P�:ԉ GBK<�����,6�������!�r{�b�;�i�����/N�!S�t�'�L��G�4ݟ}�AO�Kd:�	�aM�J�!�d�3|�Hb��r���!��=�uNe����O^������"��A��7�v�ԮG�30��t����=�
�(y+����✳��(�!�8#߬i�Z
�+�ƵOQ����I�C��y�y��N(�2�Ec$�Y����i\9n_����9�ea�^���Fz`��B��'���r�ph%�-���S(���s���9eK���n~҇�M�<|<�����}�Š�\�E�a�Q���S�d�qDB<��V�yN��l����n ��w�L�T���|��ك����@EL^�g��uE*7,�z�a����ߍ�\NNS�a	�u
IT}�ۖEL*��-�7+�ʌAv��".���2�4�hNe��;X����w_�h'��ŕJ$;�R�,����閃��m�H)}��L�mj����W��"~������K�ONGP(���Ыʑ��ڣ_8K�&��NNߑ�a���{�k]疝�؋M�u*UT��������jI�Ƌ���������,ߞe����o�Z��*�lkJ�������$�B@�Y��`���2�l�k��:��z��3�M���`0��*��G��aB>���+q}�9���d���5����)���� �I��2�$� �x�K^nw;K�˾3��� �;u=���2 ���Bo�VG�z��;Y:��@�����Xխ�����J-�#Q�nwMB�3�M�c����L��?��+�Ύ�!M�Q��]g���F�����H���MUb߻~�C��W
[��vO��|8�h"��>l�*iK=}o�][3��xՆ��c����Pt�Μ�\ ���ǟs'�R���ߙ��sH�UC��� ��G��׈���5G�3��cw� a���J7��" .:�p��kaF2�����+W�}C�L##�bW������t 抋L�F>,���A{�:@
�NF.��L�;b�WUCgtSc{���m�p����d�[(9�x�1	�B�*��+N a��|jvv{/Yg/4�Bi�P���y���| ���ݍ. �r��/kѸ�H�����u�=<�#k9�ы�����i�����x��	���y����чH�JF��GV�"�Jb:}{<�u|Hm�`�?������9�v"�5ٵW�S�����\�Q��uo���=(��I�3�o��G?$#AH������Gj��ع����%���-ċ}����b��\Q �8�:��p��!�k%��P��m|7�]i�YA�.�\�Vm�T�H=˼�@�t��(�`��*�sI?i{������C���p�W����k:C3H%b"~��&YT��z�"�`}9����!��H�fn�>��%4t�Y���H�fy��y9�w��qF/�݇`��8_E����m_%�_��ɜ�W��L#��ˮث�)1���\y�s�cA��xV��ädR.8�M�S�W,�g�07�P����X��~�Z$E�W~(����t6�00��s�N:={��WtA߽U=��a����r�#C�]�G��x:�J+�7ޠ�{?j��P�����ww�֌�n�b����K�@wk�\z��z� ��k��� �U�Rpho�k�pI�8̖]����JnzØ�}Q��:�؟sOhd�Tj�}�:��M�0���&<�g�@�m�4t�rS\4�F���V�,v��~��;���zA�>�(4[r�:�V�C�AG	�Iy	8Ń��5�(k���R�}"s�Ur�z�2�_&���@v��.q���;��0CDU2�0k�����jy��S��.Y�L�6����!�֐
��9*g\Y{[h��tT!�.�!�Gi���s9�lu_�i�KNLn��%b� ����*2�p�Խ^V|��� @����p���ʓ8e	ei�W��uD�y�Wc����ώ�SDsJ[�P��ͨ4])���:�g���[+X�A�G�j�h90}v�K�]����$��}�4�0̯�%q����PP�r [�cP8�g��1��*�E�F4K�b6"��Y��t�J�5�������ŉw�U�F{ѕ�WDHkE�%�M0rU�J�_ɏ"�¼2�-s� 	ag����V�)�塃��Gz'ru��!T�Y����dMrf�nl�ړ�2~�jA�w* �o�D�	ON���\Ɽ�A%},�NTK �(\��Ņ��M<�}��W�Ɛ_�&OJ#�ӭ��-ҝ���@��x$�$Z�5�d�3�4�_��H5��G�T'��ҋ=�M�!I��1��	!�L��2hX4���_E< c��h����_���\m�j8H�����}41@�oO䤹&#p�t�����"}^��t
l��\ɖ�a�)�=u3x#V4UZ��N�tr4W�Ƌ��L}�~���@����z�vۅJQ��+X՚���TZz�q����t䶣�
��?�xeu���Fa�rLk`�׎�0g���щm g���u��{���j3����\+�<Ե��<@p��p���nU�;w�i�"\�'�
94�$����0��8'�aʑ� ����h�CT��GU����W���\W=�f�*JX��c7#�ֳ�����S��ɱMa��̍�{��rfk�0;���^�E����NE�ay	��m�<���U �o���3��P�i)��m���0�g�\(w�s����],��&3'�:�ܻ���R����~b������+��tʼ����!S_�<`.�_�!�toő4S%�C�t7���(\�9@.�0,�'5���!�
��*�����Nflp���"{ݐ����|X�L�&��|x�c}���h�%��8���$
��c֖eM�ꄣ|��@����͋���N��"��\�%��m\�~�X4�����f�ŎE�~16b�L)�,����e�^����o�<�;������)�r��k��2�����q�1��'���Ѩ� #��d���5z���S��k-�W�D˩j������+�0��'7��\�l-���>��*E؂���P��/I���C�^�˨����'%/��Z��0�B:gO䜊�|
�_��V,���s]T�6g�G��<(����2ǂ�d�^��ٟY����CYv��a���$�H�ӎ$Ʃ�H~7��/���7�F�#N��Ϸ�����A�4�U熐c�̽�V����`]uRnxR+��N��ᄩ\��b~���(�%&H=��j��.�'��2*�' Ò�}ŮuloF�>�p�}O=����3�.�#b���g��V4zHb�5Wݧ��1qB�Y�{��P]�4j̆�/�M�\��B0"ջ�5��K�:5v�,���Ƈtk��9�x�g�[�gp�?mnLw��^�:4S�U&�"�Gx��)Sƞ��z���& �N$��'���On�������$%�����&e{L�(�nkCi�M�q�8���ѫ~$=�"f������'��w^<"M��q��>(
Ď.�y9���G�a��*�4�b�B�m���me���{���k�o	v���
��8�r}Y݄j��;m�?YLGaa(>4Z3����7#�`��+5���7�)���;enylZUY���|G���	�lIw�i�LCn��e������ؿ���&ݡ`�V���H��� K���;�IN��,m�!�@��q�D�_�X�6���_.���8̘&�Վ���;��tM$�B�Z����<[�d��m1Z�q,��)���
	�� ����i-��e�Os"mH�/��"W!�s$�d`���Y�R�J&���������ƿ
K�����S\k,`0eÂq���/rT�&;IN�e�ô�b� �����ym�h��7�_�c�
�_��w�Em
{�S5�Dn�_#�v�;�*A> 00���{�q�呅�a��k��vψy����:���Ҹ������H��� 6� �-�<$9��6��Y�k��,��=�r�\X	��g��-Ҩikd�	-�5gU96�9��:X5�]��<}�������o4��D&�׻r[����\b#���M�\RhU)���:U|�-��"v�%ue�O?��� �Q۵t�������Ǳ��h/}�v:�Fد��B���� T�B�01H��;tOu.w��J��f���H0���y��(��V!��rwY��.�H�A)+l�u��~2���^8I�ou�KyMm��9�+���>�BDQH�]�g�(� ~�0���?��E@����K��Q��Q�����>7wl��`���`'\X}7L��]�����.Yh}㙀T�M���n� �o4�E�ˢ��S�ʿ�_I����>Ŵ8�>�Ix�Ų�r�5��|jC[(C����''n�*����,�tF4L��$۬?ݮ�"�<�F���0}�!�o9�sC(-�檖�!��9Fb��}
�29��+=�����ùE2ʄ�0�t�����Н;����뚬O.�8���R��zˡӊ�����(���D#}ֻ.���y����z��t���p5�����%��W`�߃�>{w`%�,�evS���Љz߯���ڭ"tE����+ҝS�����i�s:�pl���\�o�R[�	�@��L�҄x��+��k�M�L6h+ב'�w4�4H7Bl�eh%�[Ҳ�*5���%q�ob��^�����Bq�x�챃ńܓ�ځT���ԏz��fey?[)�YG�����N������E����6g����MYO��~R3��?��B����ƾ��gX�Ķp�{#�j�b�4
�I`}�u�~�=~栎�T}��E٧e`ч�M��K|	�t�Y5�:�`���n,�T$p�%' ��`o9cm9v�"�y$��W1�3 ����%+�q,�������h�2�,� m���(�[d�`/��P�p�{兰�kѭ�C/- '�r8�$x���w��'<���S���I��G=��a��_�T����<�rB���&�����5���{'L�3����y�s`�͵�D[��Nh���Z�Ryu?(b2P�gYtn�XMm�HQ�T�sHq��-�pe��7�*��ݐfuK�@N͇/�LEֵ�X����Ċ�h�#�O�ڳ.��>Z̪����J��53||�(��m�����X��~e�3&�.V�Ax����Θ:�y��
h�L��^�+gh� q��
��
�g9컩g�_�G*\k-��C
��g��K����` ���Ё�؁���1S��^�X� ��`�Vg���!�?e�Br�����\7����3�f���_J��/ҟ:i�z/^RG�7����KJ6�id�h�7�y.f)m"�"O�����q���X��LE�0��?�^���V��<��ቐ�	�����
������2a�~=�4�O�r[�G]�Sբ}Q��ߨ��	��}Д���4ZC6 >�tm��"�����D��	����̲�h�l����&�i�����q�$ˠ� /�� �Fq���e��$V��_�)�g��Hpt��
�2<�Ș�HT��@����S�/��+D�j�h�?A@�(�xL�t\bZ7A�H�R{_�KӲ�������E���3�mN`X���ZL׵=�����D~�p�TW"�-�6�����]s#�uh��(�'M$�|��3,0jc�B�kC�?>��)�x�T�£&��];�jnA��d9�~4�C����0����&�n)�i��#,i
����*��ec���5����q��-!��Wf�F��C���VҒ����Xf��8������> �����m�B�bi���s6����_G(���c���$Rp�����*����^�Ȃ�W�j}�����qT�F`\o�}�eؒi+��`W��VW9��yѾ��������^E��oy�2�Eqc۾A�����AxB̆g,Ѵ3�#�*��U�D��ʛ;�o ?�-�J�h%�U�z�@V�+��t�!���~�]䝍�1�2���!Ѷ�M�Y��g�w9S��D��u�߮�d��iAE��h����ξ��]��f�"�񴀨��8�Z�S�Qތ��k�������|G���8���ld�����S�'������i��j������Y9�%�XlxVHYEB    6184     f80W�\�ds<�	���/��H��IC�"-UIF��Z�G�ޕ���w�=� �(�������X����D���Ls/�2|�|V��H
f[��;�" ڇ�ܫ���^x��\4*d3K0��!� � ������Ze>;�����]�O|�兣f�i�D2�l����~�.���n���f3Ih�S��T���ё,�c���ZPZi�*9����t�����oW�m@z�5���0&B8n#_"r�D�.w���U%'`av���sU>DHC��h*������߷�6L��+���"�� �\�|�wW�Z�s��{�K�ͻh����~͚�
=�[�0��XL����N)�\>�>u����^�m��$�Y���=�o�������O�%�T�D�E��-�/cL������|�������B���)����ɟ����~=�q�Ŋ$���:#���w�5��}u0�m8I��fp�������ܲ��,��l+�8Uσ�1������(����h0h��$X�.W��Z]��|_���B��X�A��#��Z�['��P���ׅ8[u��r7���&Υ��,��/������ ��ݸ\w��G�r$H�"@P��l��j�|�ނ�4&ǌ�;�~}��Φ�U���͕	��z)����� ���3�А�)F�ǔ`���Ɩ�f�Sm�8~.(�P���A�[ɻxd�:߸a� ��L�I�Ā\�z�a�V�K*Y|݊U }͸p�  ��
q|�ξ�����I�f�h��ڧm^���o�F�`-2�e�����u�_OAR��)S{��`�%��Z��ԶM������9�_���u�����bK2���u��5k�����w�0����]�U`�{r�uP����LV;MyL�j�_�Ǎ��x!!����h����jL�ޘ����c��ݾ�h+���$�Ǣb�9�HX/1����;���X-�%Q�YTx
5t� 0^���Jց@�2ܱY����[t벣]�B�:ʾ:mE1���#���I���T˝�,rO-5�8��T��'�/�H&�}����sg�Kr6���e)F�����G���n�l*�9V
R�^���Y�>B*/،R�K>y0PP�6u�s;ݓ��ck"�x�V\���6�vܘ2�^s��7(z?���.��ͱ�5�P[l8�$P��RC�5YCe����5����V_¼����'C�:��F:ؼ�XS���V�a��8�%��z��ǎ����~8_�&�*q�?���D�V�t;��yT5=��G�������@�5=ƒ��8�ё{�(g(��
I��~G�4q���P���]mI͋�&���H��W:��~�=gIM��XJl����h��ъ����.s|�@y�ageY/�7?_bV���={;�#��1�9	)ނ8��au)���M��-���z�/�*��b��!����]b|V�NZ���j>�ø�$�2�Z��5�Y�m=Ҍu��8-;�?�y����>����Y��>�7�x"���Z/�����yƦ+�����)U���Zm�c��\��L�yQ1��ً�'R{]�]��ht�-.;&ރ����l�$�b�~��m�F�+Y?��Mz�a�F����H{�uݑ��� �ìTWL-D������[7�n�W��ܳ�E����J��3t㜱`ǀ��[M��	� �µ4 �G-�K�c�p�K����a�W�-R��s��c�h���,S�ĩY�%���yf�<�_͆p���b������e��N��2³�"BC��k�W�gg�	;M���V� �JQe��>wJK��~^*d�g�����)r�A8Y�{�t��	7���s���V��Z{ϓn��� ����$���{:�(M�"A������� ���fb��k���G!'ꁎ�݆QGA��1�B�1��Y$�3w�f��D4�ꁫr�6z��������ͯ;���464�	CO1��1��"�o�ؽ���(��rKnh0�=�/�E�ѹ�10��
��7��w����kf`ݺ�11��y�cܺwWG��P�ftg��[v*�_��jd,e�"���,��@ �P��6	 i-f���3� ��!�Z�tN�-�|H����=�8��1��/A��.r����� NQ`��]b�^�����؃h�onks��E�"3�}9v"��4x�)i��l{�}e_�Q�V��a!Jw?�5||�8�����P7�Vw�'�*��Q*8r3E|%i7�ey�RL�\���*�ܷ)K��m�t6^<��M��$p�x�p�g`���iG�۲�e�R�F����Qm��9�g�����;��@;�����ߵrJ��_�ucz�i�-��y��h��;�|��S��Oa�(~e��?�|}��(S�tqxtgΉ�ʹ�n�ttG�� 4I��+ԭ���cw�~�F�}d�\C�7���F���CB�u�R.m�^J~�P�ˤ6du����|c/8����嘬C�;���/%���6v�^ �TZC��w��{]\�_�f�=ޏ���O���Z/&�mj���QX4[��;"��f���-�t�;9e�_���n�ᆚ#��2�DA��/��Q�'���K���1Jy�Rfv�͚���e"I� �z�b1��#P�B��]��|-�&�9^N�ɞDvD��F�.l��B�>�]O��nt����u����ߏo�����ghn��J����c�x$zpx������/��4h�~��J�r?1��%h�n��I��O���uT\�.#	w�x�V�{���d�,SPU��y۽iry���W�4������t�P���thпW��!ܞ{q�<������u�Hf)~�o)�Ӯ\䵂LNO���bn��]r�y��������()�1�#]�e�j�]Z�D�\�?Z���y����BtOf��Y��B 8�u� �6�q�Rt���B�f�]�3���|3b���ﲧ��B�3[�� a��P�I�Ŭ��3!5$�<�pl�}t�cP�qqw��7�p��E�w3p����r���&cA_Eܧ_w)sf�Z�DD�ק`�SprW�e�"~?��IJ���;+�������bJ��6�])_�cW�c���~��i��C6�"��#K�?f�E!�$�n��m�Sc>�&8u���^��y[�����!8�!�闸?%��J��^(] ���u�S��Vv���V*k%=���J�W;E���n,�Uq%�Gj�|5��ºk���@+��9K~�O�e�z`����h�?j�[~o:to�M-�_XB2l��f�*#Q9<��� �yQߖdұ�a�h��6	���2�5��V��4	ē�p\�P�ze��w��}<������*p惛Ҍ` L:�7�">�oy���I*��"��S��*�0 ����L*� vǶr��:Hg�\/X������n���ɍ%���W	䮨�q�)�E��l�E�r�N���A��pu�>Py��}��2v�_�DO�nmA7���y�?T�;�]��EWG-S5N��B����c���n5>b��T2���zJ�|?W!���h̩O��-����WN�Q�C���;�G�e�g��Yh�Wlo
c>m��A�%����4���SW��������V4�K�d>��7�ǈh�K ����5�ղc��N�P77�>� k	����i"Q�)c��5����|A+9^;���$���x�0�֘S�T�'��bPB�����7��֒�o�VLE]��b���x�\Dl�8��>�5]���ơ�>���!A����7d��׏��]
�����vR�L:!�4Qnʥ���vY�Z�������b�	���N��UևEr����_��â�<�3��;�d ��qD�T�~X]2 �g���-,N��