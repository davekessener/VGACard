XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!{�!K�kb��)K����a��ҽ�E�Cx�m3�����N��F�jU泰��}|����F����쵉r�]�wV�
�,2��8?-�	�EL$EtW��sI�LX����3u�r�O��99qf�n6�U�/����2�0��T���&7�k����8��ַa�^�{�Ʉ��O�5=A$��%»V���D=�mO8�}*�'S��l�g�e�v��g�|�Y��h"j�^P�b>y�$-�ޢ�R���I�a^цL��\��;%��u�g��9ԟ�$J��aݏ����R��)�/�&��V�F7KvPBZ�6�J@�wE��R�ŧ8�a��O�#/bBZJX�T^9���+1��.ߏ�B�5�����x��x�.�"k���H�'^B���x�Nl���<"1N ����f̣q]��E;��y(���c�K�ԩ��/4`z�7�&P�M���T#:�^�|s��p�rZA�s_0���P�9�Y��?��ΡU�"����"��N�O����6V�9�����}E����t���ӗ]
L�h�>RJ���M����8�OC�AklM,�k"�3��A����&���;���Z��ղ���l�_'f�6���u�f�B��3�Id7�b=˽���+e��j�3_?���V�<�IC-
!��n L�m�3|ȝ��q �Dfۅ�[�!�R��bl��㍱f{��0�xĥӇ���:���p�kk�����঱�JŃ��++�W?�g|�Ƹf��=�Y�X��	+�[]�
7�F�2@a�\�X��XlxVHYEB    fa00    1fd0�4Pe�G�He���0��b|q΀\-4���G�r����������*�j$�3Z�������]
[��S���X�|!蓣��G1�R�z�T:] q1M��do�?���Qx�f[�Џ�.8�'�e4Di�ېz�����R��K��v��(�+6�c5�`m/�@��`8t��2l�lf��Ef��Q��eţ|�xh��Id���T���!�UUj�lŻ#��p���a/0t�X���ڛ��8����(~�HW&�n|�P������"Eʱ��G2�����<̦B|�Q���a�t�g쩔.8�$���C���E��V;O�Ħ|$(�S��,��!�)AN��YPG��:��a�v�u�+L�#�K�ŧq���=TB66��IּR�%�Q g<He3��I}�A)D۹�4�{��˷b�j�Y����,��k8̄	�JX��0�i��[[�,��@�H���RƎ�bFs0�dy�(kg	��eg9��w�����,g�#��@nry&? �q$������;���,yD��o�{r�����V�Q_�`s��\�p�Q���,��u���)�0�`�9�T��%��f�OwK�W)M����g�C'¬{�=�)�.��t2��"���~���b�>�I&Ik~� #��Y�`�NH���;p�9�� uĭ*�2�(�Sň����8�H�x�6�?� 9����'p�5O����p����e�
O�y��)U�D:�kw�����vRӋ�K'������7�+\K���_`<+$85�c�e��0�c�n�K�4�`J@	}��<}�_�e�R�BWL����G�0v�P�5�,����"�@�,]b	��8}�f�򍛟e�ә�o����t�`��ˇ�#��3�?��g�o�q�"is��=�D�޷b�e�;R�m�N�m��p+��2��|g��Ѥ��b�+Ij�"�<ma��_8=�������7G�zuF�]KVR�������!"z8�U|����jT�BG�S�L�Y�m����0��	�x�`
䋊V�0� �QSt[�0_}�Za�Pcъ1�g����.��%~�Y����B�Y��O����Ʋ��#Y���?0]�T�a@#�<����G�H��c�-��3ҥpw\(��Ĺ�}��4�Y�3���`PC��tS�E���`����b\�'�'���z悓-���/�ȕ��	���y��n�� ��T />�:K��qo,ZI)�z��]6A��耛IG��U��h7��R@�ʅ�߁��X^A���d�Nİ�T���{�_߉�\!��C?�t-�O��b�1/�?7_1C�ː ���έ����?��(7)ƥʏ�^{x�[�G�P/*�����xף5���,e��8��u`zl9չuf��߀<����5��z�J��W-��K)c�cU�gH3Z&$�k��\�/�d�L�_v�e�V	��v������\�5���tT�����D�s����޸r��n!�C�g�Tu!Ԇ�c?>�C��w�ۋ �v����t���y������ �
�D�����@�|�"c�(i>�z����nl"H��};�`ʳ6��+S<B��4Μ[�,7Zmӯ�Lo���@���.�R�Fĳ����/pY�0���˒�I�&A�I���W�N�@7�5rC��R�H��޵@�vX\��BS�������
�3���q<�0�V�"e�ï�Z��2�J?�A��Ó�1�N*�]z�������+�6���7����{�_E�[+�g�_8m�J�\Y�HT�T6.�o��"���?~Ml��:@��Q_�8���
7:S�ߓ�)��d��sLÀՠ�s�BL�S�À��s��r:�;M���r�1�&RAB$P ���:�K�r���s�璸e���@��2tz�}�����pA��"!��Q�<Y,��X���`����2��ӕ��_���Ʋ�zםJPPѧ�k)No1�]p��t]��`bx0�~Qʇ $mT|w�Q=��u.x�O���!VR}��p�t���	>>���|� "��C=dUgh�]r��qǶHр������L(j�d�Xq�Ͼ�����]r�$��(t���e�{4�{{((�j}���8���Ζq/�5�q�. -n�r�9 ���uQ&�F�{`�y�4Ɋ%�/��\J~���.L�k�|��E.�m�{Hvy����'Ѯ��!g�rC�*ȿ�L��~C#m�ǂ�N�=9���8�h0��jMy��TZ�\�H�6j�,�Wy���\a/fj�w�i6��t�1��V�0�Ħ�d��갘T��2<�jXKy?!64��8+脃�XB�K����xV�K�L�/j�Qp$Xj��x�i�a9F����i1������@o��Nvb.�v����cS15��?R�k̶�����k?B6B,����-@�F>Aϛ���k��7�j��W������y�Qw+�Z�r��Z�6g�V�B�au�uwe��P�$��C���������`�y^�]��4ҽ��ɔֲ�b+��
�@��L���}6�^�$X����@�+��%ᘋ�3�=��4w� X�ג<ۇ����Z���b�1zp�E��e4��Ƴ�2�X��r=�O�:biPzC�'#2RD����}IoX�0c���M?�K�l��jYUR����[�VS�M����O�$�*����(E��	.�.3w4r��	
�"�R-��b�5���&���m��)VW�zs�*IxD�����Z!p)\P´,��J�ؔ�?�zm�M+<@�p7���a\jf�K�r^�^��Ezm�p��`�8#!¦lQ�0��b���'m����õ�vG{�`��x@,8���)0��C��-�Ԭ�H]@��x�V��:-����9VBSR	�+v�-���\�$!\Z=,���c�\�d����̚қ�)��^.��ڭ� �j�n~�(24�zu2<P,4T�ߤ�e�Y2��M�B9�(���� %Ԏ<M?�B����k�v��V�%@r��seq3m��֋N'�8S��0Z�V�Y���n����{�qa",í�Ogr6�b�frك9�p��-q�"��z���x��!�7UC}"٣ �]�|ZG�Nf&I��|2'
��[-��	�-05|����f�G��!CX|��Xz��M�j�����(5@�M8�Ӥ�5"~�O�Rm=��{sFp;�����>�PJ�QB��|@�鉿.��w2��	�@ ʥ6*������M����� ,_`��p��}�._w]2���x�eZ�|sS�9��<�^H�V���jhS4�/ɺ�`:']�d��;�Ӕ��Ԗxk�̄P�s1�	�#٩��	�w犎�f�[�E���_�/��e�Sm*I��+�������r��|؀����,|�(���vY�j^��+}{��0羊��u������^F��	�����͍9ɒDdn(:r���jOIwGtg���3�rt�x2�O�����9rWF�ѣ���bQ@�[ֆ�ѻ�r�0�ig���N�}Ԯ����5����`e����LlMP�.1���y{�,�:�^6��\#�� �3r���a{W�r��ש�k}��]9���N�u�"�`%��>uB�`����l���ZÒ�jr�$#�Dǻ0��Rlˉ��O���F��`Tڕ}G�a�L�'���f��J�����']!K��ހ�����goZ1��C:N*��׬�g[~y�g�3�h���/�v�����JM{��q�~
�����8M�{k��(�*E��"�{;�����H=���R,v ��٣f�-`�]���Es�U��t���ӻ�w��)��5P�[�߉9Qg���~o�c���]�&�K����_{�Bw���Ai��k��!���鏙Tyt��W˃�>6����#����E�T��>�u �(��sU��I����� ��}[J+)Jv�����.���s�m���5̜u$�y%R!|SIz�F��(CW�)��U��[��J����S�C�{=.k��؛_�$c
V:/�kK�J������_�����rdS�u����M�?������yd1��� [�֛D��4�� l���fZ��m��l��pE��g}�:1%�:!�e'Ƀɵ�Ñ	1SDx#���w�й�ȼ<�h�]án�����LK/#�0��guhZ���me!�9�4��'=z֎�w�EeE/�?�k�/�1�gA�M��[]�Z�ޣPbx�1���GS�*8�|x�jta*�h�Ў���;c!l�
�C���7�M��`D��� ���^���.^�W���"n�⫝̸��.�ց��D�@V��O�LԌ�oM�{��>�{?T���h��I����9b>1K䤛�#3QAO�_�E����иQA6�� �=<���k^@0��k����ĩ�i�U	�� ];.e
+��{�u�����k���Bl�ks������閻6��F(�\��p��;`��|���_ƍ:E�I.\���a6���HP��c��2H�hzq���{�f�j^�c�hh#�lԍ���k���K!��bG�v�e��2����$W�iX�r��_I&�78Rv��A\�[Jv��:�B�f���c{V�~6�?b%�.P$_��ѫ���/����p�ZFQ�]�=i�U���b��dhP��
GS��ŽTu�1��������i�s%Rѐ7�w�`�L�Vqc-b��N���*5?�-���U���
ó�\h�mҕF����ܘ���앻�U~@s=%� �){��0VS�L>���ݦ�e�9�껱`��T):C������|�G�[�}{�wO�A"�B>��1)]����/TO7�V�?#�ٓ`V��p�J3S��xC�&9�x��3U_�=������%q�ze��M-T���^1����u/:�p@����ѳ�w�t踾��w�\
�������/������pw����$�d�-Zwꄸ����R���H*�������G+��u4g`�7G�����;'�W����(���%��rb�t�Hi$żr����C��E��tyĈ,%T�V�D�ꘒ��i}T�I�P]�;I~�J�m�c���/��H�Bd��-Ul� q6�[�� >p�'g���ڙL�q�skT���] ���b�1ăLy6��>�e�v;[�f���#�皺��N0�Gg���e�7w�q"a��ݺT�5��摊.�^mo|>�XT���L����ݾPR�i�R)�T*��� <%&��`�?�����@�6Ӵ��T��*Xq����֛�`������.1CH�d|/X��B�7��'#��:u����iRh_	�{t*%/?�vTS:��V����ҭ	���6��q:Oa��^�vaĖQ���G���i��A~�4gǥ\�H��9/�A�K��ӎ�L6v�t�[/�s8׏��V;Ͼ%��v�)'��wcҳ(g�{i�ˡ�W&g*�|)�o �fU�~��G�Ȏ������"%9�p^�t|�i�D�۟Θ���h̪W}��+��R)p�N���&�׼X{H#u*�<1�v@f�5<�iA����R�CvG+��� �}\Ϋ�y��?�
�-ɸ�\%޷V�o��n �*���T�n��GGT��~BY�@�<�N�`�[Go�����˛��VSh�/��;�!>J�=w>��[-�?u�~��0�ڇ%=t?6?��Q�����$��L�2�<��xeETI"d�@L�����}w�d[��M	�����@k ��4/�����UMtꕅ:�p��3Y%���{�I�� �#ٹ��8�_
D�������*!$����-#`Yq2��\l�1�tp��8��� ?���t/~Mp�B$���� B<:��7��3�s�x�
��'��0=��}3�-Mo��u_�}��o����-��6�gR���	7���F�ܳ��碢���>��������7�!EP����+,��������|�����}�__:T
�}���qJ*��4��L���	G;$���(�E�{���A��v��n�(�u"9�I�ZZ3Sg#t��Y�*ѴCN��=x�6Qh#��j'���V�������\X�f0G达�V/�-M9�^z&��NOs\�P��1�]�`���C �$�ݦ(�L��l?�W꼹������h��c�����^��D;��~���D�;���򃟝�ǭ��h:}"n��ہvEp^֜�z�>��-6��r�d��S�*�����Bq�0+5Y\/��$@�Ŷ��hx�T���$��R�)�6S��!� ٿ�B
�'6���P��>Gm�*��~�X��E
��gj��.H��o&��`�S�¥/�I���	��!N���M�~��<�u�1F��쩁��>Œ��������f PD0���ڋ�c�������$~ � U*z�<�
��uw!Q�"��h�hY���r��$�-Y�|�Hd��\n�)գ�n"� ��vL�ҝk,�YI�f@g����{E���ۊ�X\W4��Ҫ����� ��{�6���G��#�����$~|u,��0ƍ�����	}�IH���#2zd�N�͔�,Q�	�#����Z4�:�ʇ�B����Sf-I���Nm��̔���MYl3�倏 ��9�'��
Dg9��Ǡ�� @�E�V/��#���|x]
�;�������͵�e��N��L�������0�,�Y��2�>��u]�����H����!H�߻�Fq�uf��q��- G2�λ	'=�^�K�g��fďC�S\p���9x���Gi
�J�`f����J;�.�JQ�M�ݐ�M��?<k|W 8�kRO$�4����Fצ���3�~��Q[�����%9��R?K��xɃ$ �a!gW�������[l	�`�|Ğj��e�ΰ��������N��:U�f�I�/�UX�T�p��l��Kn��'�os�&ʚ��pE�C��<���C�J?m�l���D�lO�:�X�u]{���T��?l��dK��G�1��0� �&Ήt�k�XlCr�������}�S>�F{bs��,�`nP)���p4��c����e��,��ߒ)�5�F>_��m�H���ۑl���ڮ���_�J�w��I�0�<�:��g �'q��^2��f�H�Cao&�̹M|�	��ڶNz�0�D�k�f�cF�����	���ڤ�ͰFg^�N�qM���/�	\�u2gXh�k~|�W�w�,���T�/���	�TIE6�/r}��mD-���6A�察���49�^JN/p<y'�6���z��­+�O�d߈}E����F ��q�����S�rB ����ݕn���h��Il�3W�Ԟ��tʭ	�FL�l��έn�M�\��:	8�O.�ǿdLX�ȍ��{��\�m ��.��n%�bB�߹C��	'+n0i������k���c_���b�a�G��S~�܈�s��6���wm4G.[�l��o8*���]�T�\aLk��ƿ�"�h�jO,��BXh!��.6%��D���YM��e�
L�r3�gy��Z� ĭG�Y|�
wPߚ4ԏ#3?9�NE�Z�D����`��C�B*�K^�ڿ���~({�"c�\�҇��v甠�Cz -�豦�k�:�_�D��
+�R����m����ȍ��D�ͱ�*�f�j`|�� � ?`�|BP�p��� NWل�%y��"$����q�g}"���q���D�6�P���܈�q���%��^?�h�fN�yf�|���E���'�����W������%{�����Xf�`�[�6P;��?��q�,�8*A�D���ʅ�mEk~��5B���F}�d���&��Ԕ�WS�x�_<���*Lt.�9|lA"��_o)p�#�3���`ឿ��&v�aV�w�.�DVյoR�є��A�z[�3�����Or�gO#�FM	9���+U`U;���LiF�rÃ�`��k�4&wl$�G����G\$�E7p�1At��Ƈ0�7E�~�<L9�y��;�H���9������7�2d��H9���=�XlxVHYEB    fa00    1340N�B�s�i�9#���5��!X�/���}д&Pd���T�V/�T�e4�p���ʸfz�=M��ݺ|�� .K�s�-�>��ui8�wB���ח5�<���Y��Ҋ4��[p=pʹ1�J௑[gY2j���>��i��t	L��œ�Ҹ�'�`���NM�U�.�]�y��#d��;j��N�h%���+������:f�)�v�Y7p�i:@bSD�@�'�0��%O �]O��?=�6��zUhB��o�N���twe}�?t7�XY��E�(eRpX�h��Ie�C�>@^���,�Ѣ��6����n��(j��2 �Mz�1���J��a��@���Ok�١Y�,��uU[����6Z��.�6��S%���3��o����L�;��Kt[��K5FDq���&�8X��A�Smeو,H�A�^.�_,��4��f�I�ZL�D{�V����iwR�l-?"-����&y,�C6	}��i��+R����X(�,�q9f+\�U$���:V�g�a?�,M��?U»��8��4Ȋ.Ka��r�����e;s1�Ih��Ȍ�۟ѫ{�9x:��3�K��e-������ a8�<Aw�p��$�&��Q���s�t	�G�<�A)X�����d R�0և���98�#+TGy���˭��(=���K�x�Y>�,s�p5��3٠v���RauI����a��;9|�kq�AolC�p��2�a�Ma�����|��(�~��m�R�͞Ul��w���CU��34������DPD��xu�$��(6U��`��s;[�T�^�����v˕αe¢9KJ���.�k/���_�8��N	����%�Tzz�1�.zr�-�E8#ֆ6��j��$�	q2�u�뉍]�yu5��Ėr��yq+��'�ʔdc���2�*�ICi�������d:<��v�<����zI��t7w[^����f�(,�v%*K彺��R��}�L�fX�$�һ�R�P�Xu���C��� ��<���?���W�g�] U�[�`�9��o��$�z�>MZ��P����+W��d�C�Ap�[Z��9_��GS�i�5��� ��c����-��M�
��>R�h�`�P�������j50yShcئ]��T�a���	�H�+ƐU�gv��S/��,�_��$ �>)D�;�,��T-DrIo�ٰ�n�j!2�,i�U5�^OW���F��5X�L!t�Tp���{�^|�j?"�'�{AAЃr�{�*�T��f����!��?���w���~GX��;�F�*���"t;��<���e[��Tz�w�l�quY���8\f��^
)!0L�V�M�(�\�-�p�0���1h5�u&y���Ρ��Cf�`���C�pR�I��Cs7#k�EKPn�۳��1�q ��(�.�P�̭3�4�q$���e18Ìf�P����2�Q�����Az�Ys�k�g6"���~��K!έ�o D^?�vh��)�a�	b\G��z��+t��*K�`d�̵g���6�΁�[>⥻��E��V���A�lH�[p�6����V�׃��O��H<j5�{ϗ�Ģ�h�ʭ@�A���h���HG�}��W����Ԁq�X����`敱#p�H�k�`��t�a)�	��۸j�����q|[<ɈD0|���C� ��$��[W:y��Y��Y�
��*.o轕�G���"�Ջ,�ԝmc����67;D����h��?>[��4Mߴ�eM�-7O�y=%��R�.��2}�[̪-!�!�DO ����=��C�����fR	�`�`-�F�	�]��*R���M���M� ���sp!8\.)w¡1YL�=8̴Q�)����Bm�[ʛ�U�{8����ё��f��d��r��<<tF�7QL��B|>��wk�AZ-g#<N:��vb~����~�&��w��;"��d0B|�^��z�=9�y���1�cU<{*Qs�K��D�h�8r~�vtd��_4�w��!�L��(P��r�L�\�9��wB�A��	��8�����er7��8>.^#A��"`'y�}����;|Կ�0��NrG�Gp�p�xIO�c�����ȇ���x���ry�7�\>��,R�w}bit��(�D}���zL�t�q����wI��R��o��kfcPK�oZ;���}�䲖�\�"�ԝ��дL��/$9��2B4�aPde�����1j�5]�omWR���Ipz�'���&}i�g��b!61H�o�o`X8��/dԅۃ�<��\�����9A:�u��W�BJH6�B��U�E
3N�e��t�yBu�|=��*0�a��	����H�i9�iO���M8�)��"!��r^	��� �����M??�e�լX|�1�z�<2�(���o���Y���͛���Xm�ᅱ;����2$�zew{�'�|�|�`6"]t�R2_.�𙠥e��y��ȉ]����pY	Z�����޳�:�jk>��a���$ꬴ���<s��T$U,��k�4�%K����(:%0cΆ�$��6~����v]��(̬_��g�q�U��^��O	e��[��,.�^1W�S��;��Akع�*����<���y����|s�b�x(��lDy�և�zh,�J�d/���,����?n�>���#�x�X$$��[)	��(�.(1%���%�zݾ}S*?\����G���Wb\x�X���-��C�G}o�F5��N ~׺���hy�۲��=$1��!��e[��u\�M�K��A��|��&C��ZG>!�8��^O�U�.ٺ2D�����>�Κ^}NE���F�OӍC�yAe�\7]"���Y2�ew����W�)Hx׍��{.1�bIn�����(�Wآ���s�RX���\���.�y-{�:�S��}.d����o߾�����ʶ	��Y%D�Hs�b{��$�u��&�]n~0v�c'���-Qm�H����	��i�2L���pt�o��\C�J����������ǵi]�9�#Fe��OPh�3��ia�''4@I�ۭߊe������;��"~.֍S���U��1�%)z�]��n�Q���_��,�~_�]w��]����s$ZXN�|ν)o�a`Y�!iǑC�Qr�|%�fܦ��_yꈾ����JP�����ꌚ%�w�4��OY���v:�C���}��{�=^R?}Kf5c�M�n�p&���;��I�ɽ��<0'5��iנ$��5S��Y�!\ŋ�3II������̸[K�4�~>!�N��w������^O���.���9��כ� I9��~3��`eY�p�\p8TR&Tm~��ؒ���oM�@�eK�I�vĩ���w.	�!�T��G�ӆ�KO�Z��a���z�m�U��\���c��$� ��V.&�Fz+�n�fpf�Y��5`=���l ��(O�TFk���\ݩ �J,������/[cΊ���8I��n�`�/�	:B�t"�i�ȉ����H̥��#�N���v+Z!�=#�E?C���Q����t}��!q{�^�OWP�c���y�G��"��Ʌ�]c�IS��J��L��׈p�H��ѡ6a��{��+�k��|o��X��R4bE܊V��� $5�wa���2��k^��5G����,I.��,Ť��P���p?�h�H4Ak�Co���؉Xmu����> ��������	���gh� ���><|5�$- @9�I㕪��FB���`q|uڃX!�5�F�w��*r_a��D� ���z�����Hr�通�b7k?�QN�/**4h��7u?��c�ER���4���'a������9#��2Y.\�ă��Bݧ�9�1�y���Zۆi�'���P���)�~�;���3��a�D��Y���sj�bC��u�t�y�CgBV�4l!��X�w+��>�d\ai����n�^8X��n�MO�X������x�Ѳ�p��v�d��4���4������I�D�Y�қ%Ǻ�Ć��-mh�:�>G���S��C�heA��	��{q�M�ǂ�;�]{Mp�KYn�T��R&�W�a~��j�9�@��D���Gvݶ�[���cW���i$ r)���KW�%���l^����9��9u����2�3=4�Q�F��w�(t��;T�Ǧ�|!X��x1}�e�O}N���\Rׇ��㷌��ǏQR��t:�G�6 Ɔ6P��p^�8zA�ӆ�}n�ڲ�>��1x+�!Ʀ�Mf�р�R��M�����-x�ꝶ�lT�c0 n�Vb�#��>x�Fl	d"0a�;Κ䳘l�@������~��E0�<om>�;x,E����=�A�l��L�N�)�<&ق���W�-������$	ծ��P<HUy���:M����� j��d�FP#�|�2����H)�jyL;��N����Ŧz^�����LG�	x�sKU�{J�2�,s[�Ք�Eh��ưL�+Z�V':��!S�]3�錊�ǲ*o"���Ù���D�N��E����2i��xG����~<4Ģ<1R;A���C�ݒ2'$�IN�Θ'3�?���n�Z|�[��^��.)@��Ť'8�~9�6���'����<��x�b[_���v:;�g�����g�W���Y�3��\'j�-�F�����[α��9��.H��SZ-�=�����g�T�A���@ܳ�I��C��n� �
�X�=j����7Ȥ/tܐ�`�G���Q��O�sQt\z;O�>�X�m�Q��@�X˿j�;Px���w~8L`��d~�684��0��ɎGF\��u�/�0�����9V��x.�����۵�r-�m$�u�)�W����{H�[pJU�> ;����rʒ,4�ʚ����;�XlxVHYEB      e7      a0c�B�M�d�R6���L6��^q���V��I�tw{8�#<�P��K�ЛBї��H��-/{^���D&@Ӌ�,��_��d/�9��a��~\�"qv���}���Uv6x;oh�:Vt�$Y�>�my�Æ�m��ڔ��Wk�z����_ n,�l�����}����b