XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����
^>.{;���K�:�ta�p��>�E���Ny2������h69����m9�Cg�>��L���]�m����m# K���1X�M��݌�Dڎib�S�R�ư
uŎ�0���'�X��u9�8Ⱗ$���]��+�����`�ǘ\}���.�7	���&[�g��6r��_�^����A�͛��4;:=���vԸ�ʬ杕��� D�cAб��!jZ�{;��[9NP��Nu	P,�X�*����K��tɅ,H���D8���DB��$'�4�<  F�@t�WK����kƐ>Pt= �҄@���|����ӄdvQ3�B���CN�3�.�f�!���:�|�/�}o�B����SǇ>LՌQ0�9�(v�Iz����u�tq�&��e��v�M�HY�������__:�D����V����v�߆1!��[-W0h^�:��qE ��}�N�j�x~����߳��oy��ڌtOZս�ѹ��q�w�7ɯvKL�gG߰���]��2���c}��4%�[�����c�Y����V� �Xn�͇�n�<ʩLT{�<N"����%�D���tndy���|���cE6q�����˥I�G�C���Rxk�|6��(� �*厮q �!�B)FI��\xV�D���F������~[͍W�4Qu�}z��B`��
����+���S�4�R�
'�V�@'s>�	O��N�\(f�?  �33��xtfe˚��x��KF�E�?'��M3}�������WXlxVHYEB    fa00    2470�$D��Y� �W7�W�(AM:��ME��}2�l[W�s�~� ܠH�7�Z.�E�	�a3�IjSsg�Y}��1UYo�"�r����&��[���tfB筃^w��.=�-�u�XZ���b��&�5�c��V��!-h��,�pڪ;��j¥����|j��}x(fQ��a����ѭ`�\������LC��Qr��$����|�:Zh����^9F)����H������(K�H*�A��H��+��@I�Y\�3-q��d����
�췤ˑ�'�H��j�_.�ߩ�v4^**��X0=�K�_E=#t?Y+��p��˳z���\��iN" ��Ó<觿�Ub�����b�>�����)�c�P�:���O��\�)��0�}� ���o讻6TɓL�ӰrJ��Ƞ�9M��=�M��y�м��;�J�q΢�Af��6Mu��5��"W��ԝ�hf�E��i�`t��N�V	v��x�-N-�t���H�y����l��c���N?!�&�͞8n.�������#�\�e�0��12JE�����銹G����ͺ�ϻZ��(����|���o�`ˠG\��V�pS�����[{ȦT����	��K݃yl����:�Ƞ ���^����9~�lvM��+5��8?�����јq8R�U��G�Z0ģ��+No1�&���DEo�-��G�~����|�w`ǻ�u�9��b���x�0�jv�x� ���qФ��*�m��n�A����!+�y�G��ٕ�^�	�DK)V�r�4�K8����f���JD	�2��¼�(��0�X�)�\_�Kť�&����R�xH"���"�%�J�.�Jl�'Ƥ7W]�>2V���7�iv�Y��<���V��V{~/��V��UK��`TLd�2�I�6��
��C��V伩��	����sӨ$�s��4c��&��� ��,��Ҧ|}މd�3����7̀guI3�~�b�LR��`P��h���]~�)h$�6���Ѫe�ڵ�aiěd�[� ����-�4,Yy9��*�h�֊��tW�b��mu��M/����T�n���9�єX�-��*[�E��T��I�g���$o���>}�"25��a��;Tb�.bQv}8��������Buv�+b��u��l4B�Y�Gê��"���E[���j|�P��R�<i�&��Ij���Sng�c��M>wq�@52C�2ڙ�ݏ>�����k}�o�s/�;��C��� �Wn�
cr3��g\W|�jK���/�{��'$R̴��Qr��+F��T45������m�.��Ȭ$ᑹ��"'�)��2��c)�ϔ1&R��X,�p�M�5�Aԥ'�d��R��${�i97s�^�ܤ�\��jjj"��[�35ks��:�4w�+y�M��\�Q�L%qco�[�Zw'���bP�I@��ʤ딆�&�� 30{i��I�3���M zCY4������Jo?}����M�jh�yM�:����x{O�C�%�s�J�k�� ��#=ň��� �.��k2�|�{M��@����S?DFL����'��<�{���q�{R��NH�F{׺+��`e2`��Ɍ��`��ک��j�?�[u���z?��xZ��x���H�C�.���$��;�Lfc����f.k���g��շ�w�C`�Q|E?cw;��J����8�dk�G�Ntѕ�Đ\��h����@�����5�sR%��Y����L#���f=��A ���a]Or)��ЄjT�χI��N{@e���~��-�I;�jaB�#�P��4����KأU�fP�� ��4l�X��0�-�t���_�	�"�Z�b	�*�o���9)ޟX}�eL�ۭ��aE�^�h�IQ�^_�;�ݦ�^���4��Ϸ>X�{�bw�*��B��U�0����]�N�SJ��'��#�y�>�������mi�\ ���@����Ė�q�~h�eǖA挱���%ozb�z8R�� >1r*r���ˣ�j��đӻ"��3�h�lU�q���ޕ���u��F���Ͱ��t���[1���ՆĖ�Ρ �'� A�t��3>e*6T�.N��ke?^o�0@���
l��SC�3ة+ǳ���0|ݿoPʈ����OG�=P-xR�i�$@�<eT�KRs>�j����G�����U)�#q{=�у�"v�c�k��Q��q5�,�Ť�]>u�ߖV��p"��0�g0`q������-���pہ�}�:⊄Р'3O��Vs6u�&�����}��;�qq��.�����y� �����16�J��'�H8Zd�Z�%9}%�mD�s!M�~��Dn��T�W��Ь�uLy3���:��TXt�3w"��ΆQ�[ܷ��fh��(�2"�Rm0@����g�д����������//�&-��ܺ��O���{�փW]�\?}���� �I����K=M�� ��e�(�����?�s�wy@Q��|��� �Ǵ_���0.W4��K��D�Ms|2�%�I�?��م�p@`���OL����W@cz���XJ����4WMt�z��`r�o�q\�� ��xA9,pJ�nk'�ڳ��?�۩I��V���I��zDZxPA5�@�0K��Η��yڦ���[	���VIyM�UZFy�{�;�;����^W��&��-%J�^�F��OG��R_�7��	9��~ {m�a��<v�����*����ț}r�?溥��lZ5���ͯظ����ݢ<�_-k�?(�<��CH	q���Uc���pԶ��[/�P�>Bu����5AC�xM�Lˈ�_M��F'�@�ٯP&(�*p]�E�߂	��`�M9��W%z�N��:�0�����ݍ�թ6���&��Pk�=�3l��Y��nT#�V7��ýe�R�N!���e��k'�,w�1���=u��8��R'�j��ɀ,w4��)օ4�h����v�q5'uR7��:q�@�/��:Z�`��r��{���$1i�.��G)����$��Sy�:�� ��|ư�a����ް��6.�E��*H�71f�	���kQ��b����)h��(E�W���ܚv@�o�v�!���ՠ݂ e�1��N����di���7#�ni�7LX��4�a=';4l9I�W]�Y�(�)\�L��dY�j��D=��<��F�7K��B�;Lu]C���{�ۢ�ϟ�ET����D9X]==|��#��Q���bo���F�,��vҔ�g���:���i��-}�G�P��c�q��ґ�/Bx��Ѵ��ݬ0y�a��>���nߞ�*����>HG mC��I��=���G1Ʀ/Ս�Gp44�s2m�4��0��>�X�f("�.���=�:v�M>l�e~@AL����T�7p�u�|? �2���!��x�j���ƃ�tx���4Q�x��|W�7�l����`�C�cESB*T��a� ���ש;0���#P{}����t;�QX�	.��:LH��F�#��<E�A��qI�g��C�,.�?c�k����4}��p>��<�ȼ�
����;06�*Ұ��xLDdX�Ã���!�+;ˏ�}X��pw]w69ᬧ����k�L�Z����N	�f'N=�_ҿ���q�=4��y)�q��zR8
�MZ@���˚�.�.b�z���>�����h���w��#���u�]�SEE���B���
=�3��d7B�R��A��(A !��>�u�)����e2[���`271��;��1�ޫy1�{�~�����.��,3͉mM䋏G���ΪQ]��W��;;h��pt�j���Kt�U@��sQ;�-Xv]����}�6]'� �"	�pU����r��8��;�Δ0y�r�~_�`�Y=�!��ѡ����E�U�j�l�uS�[!<#�d�V�O4�[v�]�F�h�i�[P����ٿlUؿ�@�X_���A����:erIc�T@e"j�����hQhzx/�l�!K�`���sF�I%,���m/����þ�� ��a�����XN=�?p�X1/�/��`�D=ʬL��g�]΢`�c!+P
���ђ���55�5��.�@�V&	���d]�����Mr3ڝ����j����~1a1��wU}�i �V T[��.+����Vb���$�7��R��g�A��1����q�C��)�ɗ�����y��Nk��\���aX��'4�l�*�L
���)NAXf��n��0�K�')v�_n^�g�A5�t�a*�̬�ꨤ���r�]s%��/*��c�=&a%lx.TT��3���Q�L�>�D#+57�H���3~�z}f�2l���r��#DǨ�������*N2zU�ו�f/�Yݭ�ؙ�l�nc�<��dK)�Z���i���E�) Y�}�e9�I譬��J�=�>�ͤ���fU�-���.B��dQ���]��VI�B��Oõoi��=�T�������2��Ř�#x�Q��Kb��c��}j=����y�%�ٚ���Zb�a�5�Y�SCln'gA���M�R:V�#�,h!%�Xz���5f	Ȧs^ȿC|�.)�dṒ �ˍ˿��"GAM��^�Y�8 �_���Ds	�.�����Y����R�.��9ڿV)�@�#����P�"V͆��3��������<��$�r�;�����P'���������)�n�El�Y
�DE���Yu0/Q�7�c$8R'��	��'{�[�,�%�-t^Ud�#�ՅZ�6��Lͤ�j�lG�"y�����n%T��W��
�3ì� ѫ�M���
�<��K���̣d	��{���f��t���HX��#�v}�;tp���� ���+��S<�~A{E|n|*W��'��bɭמ����v<	���&��[]A�I�`�(���Oi��)��!C��������I���������Oy�s�t$�;g3Iy�#���wD����=�<��1��av��̳��G&iօ������Ĕ�V��k�0nv�	�~Γq�{�����aq#���.�{ �_�r�p�HM��}�fX4��j��	�{t��-E<kʥgu�	�"7�I^e�YB��D\��8�sF���jԇ�t>�����Ht�F���3W�N���Rp�Y�!���6t#k>�vpD|���;Y�`�	h��u0TBB�����D�g!ǧ��#�l��N���:m)��(��.	n�n��~�;��Q]x�2|o��p�.�۳�W�����ݽ%⑐`B��q� *W��{��*�D#�3=�r���2Ɲ��^��o���7 �O|o���6g��,Yɓ��4��o]E�����+*��8���O_��&�X#/$`���[�~?Ic�xvV��+'u�Ė̵{�;�m�$��P��[ӄ�x˗J(Vn����2��#s/���G�qＢk��&)zL)!=���G��F)�q*j���t�j��kx�H!^0��v�LV��=*��faj�G�D�j旴Hq�j<쩗�ƃC	�0�\�k�<r)U.���T�K�KmwJ��S+ն|y���W9�����;X���j$oҠ�C�j�"Vi���
�5�)���v�.����P�a)�hx��,�����yt)�Z<��ks��ډۗ~ȴ���C�~yF4����n�91I����䲦-�t�9}�o&6�k�|(��4�J0������j��#ҏz���1�q|H����h��rS|�"܍�����Fb_4;���ے�43 U#L{�D��#]��&�@`��?R
����������x�8�������I���?��ʾ��(U���T��l^�0��N\�����C&�X`;�4XL�B=yE�����쬉�j��wfoW&��'��l��C�G��Z���=�T��r@���ݫ���3�l��-7~�cO��lM��lmF��
r����3��[�u;ˊ�8u~�Y��Ɵ��qш)c���?��c-�#�v�P�39�]b*G��#���爵��E'7���j�"O�J&@�i���,mW�4�-�IU�KO��j�ΥLS�ړ�xk'�d� 2�Џ	�9T��]�릘��k2l�e+S�7t
�4ކ^��@�E��&~���
���w�q�$	@��
/��k۷���sֹ'���l�鹹)4���KȊD��B�6&�֥��ޔ��W��1��gY\	U���{K�Ɩ��ͭr��AI�X�p�]r�ot�QlE�b�a��X�r����kF�<�=;�ʖX ��C���m�Uҿ�%��J�c�I$��� � �$�D�?p�?�Qo�f���G�Jd,ӜGĤƪ��*�U=�|���ZC	��<0�Q�Z�S�(GL��v/�P.&�&:��:�,��er*)51kh&�K2>Ж�bK�c9.Խ��9{��Â����Mӑ�mD)�]��.�߃�']O#'!����ȽP�X)�6 � ��F�H-�f�M�@��.�������3 �q���3o�+v` A�]��&�1���kR9�v����<m$�Xy?���K�WR������!���6��i�)_%�3�*w��qE����|�3�[��N"�g� 3U��0���W��z�C�QL�}�	-��1
eZUؙ��/0ZR��;�7CPKI;�V߰&��7�&SH�?Rw��B�N��jf��-m5(yU�
�>[�GiW#�߹c�hq���8��~,OJB��sۥ5��݇R��,�E������y�H�a�ޭx���f�U'�<�.ӭ��R/�\��h\PZ�O�d:۬�����;��b���0͂�@��d����X��������nG��|��,�����;�_�J�8m�Q:
��N{����#��㦇W��wl�z�,��k�� �k����,���(�������هǉ�����a��sKw���/���pWc�B�^)�u���[���G�P?&�x|k����!��~J�}��4 ��S(C��ʆc��cW���x�Dk$9�̕�c:��,(���{�i���~�^�H��<l_��\��h�Z6ķ{�2�j�:��h�yt�}�&�D࢝��IdS��(����j�� �!!���>rG���ꞣ#�3Rδ�_�j�� %r `4� ��^<�R,�Ej��:�P�e8>�#�I�vi�?�K����J�(��6|/���qH*���}�meᅌ<��E�ci_)$ſ�J��)}f<�6���@ ���~�i���t�z���k)(o`}��h��'���k��j"Զ؋>�!(y�R��.��1�j4ߖ8φ,�� �Mm��]�75�S���w�� �G%��)'�P����@f#��8-�Q�4�h�mƳ]Drd��5F=���x�.�D�0g&Jl�B`u�W����am������"�8�r'���]�U�3 �M��j۲�Tm��_ �mt3q�Fh�@�a�c���w�����8�M���]���M�@0-�ȧ!�Yc����YJt5��![a��]��K)p7�r���)��\��ؤ�#lڨ 5��t@�7V�YH?��
l`�ڡ�-/��-Á:IF*8yi^1���ܽ�D ��N�eW�m�tZ�1L��83������/�����߸�@\):�����?�y���2������)0�R�$� �qf�mIb���F�&�H�{������\�O_�&4�������DY�խ�/iJv֥�S��M@b*��9��8iW�>�s�y�6\LH�axJ��1�-2��=ٛ�����g$��)V>���\����̷�LY���.���mN=��cm�H�F�\���c��ybܾ�v�g�~���a�s�����6��B��/�����	Z1�k��ʶsg��
�}ï���	�_1��#�v"ZZv����in�͏����U�-{F�AEW�sJ��2K
h�ݑ�$�yK>���C����"(�6j��xjF��Z���X��K_	�fC3�DM��z"�АJO`λ]���AuFT�������K��q���-���$���ԗ�S�M��y��"� :,��e˧P�-�\i����;d7;��2K��ō����V^��Y�ހ\0!Y�a�Ls�N���$�2�B���M�����I.���m"/�E�f�h��+EC�B�����L!0�	�3f�CTJmS��c")<^zQ��V�V�.���+�99X
.�|�!��Q  �zK'y��:�ˡ$;�LDi��kla�Y�iSG~���������$�y�f��,�Z�5x�lN$�����R�fpfhg<��~1���J+hڜunι"pb�;�+�k�t��Jtb�Ө�����A�����'{������kG�K�gD.�����������]�:�E�"�k�B���wMv��XU��85�c:�=HfCU�R��W�	96�ϠVyQ���7n��8���j��4@v��r}\���+��Ϸal����	�T_<����a*Eb��݀o�(-`ՒG���6J�ep�s���6�]f����5�z!<��������÷�@�nҨ�-ptP.�s���}D�O���q��"V�]��*�ό��� ��܊m��({����2�^������i��-$(!�$8�kÄ�F(^����Po#�|���J}�o ��uA_(������cg����]��9R�V�2��ˋ>�3Z� �$��@�U�-��B�w�����G����@$~�A�_�,����s����4��M�U��^�����=�~���S�v�jZ��VgS���v@��q�k�`G�﹃�RAh7KG��16�dx���� &�i�2Ec�}ʥ�oVf�!"?�OLF6о�h_��ㅽ��7���G��$�@�zk��W�sy��������?��|#{'Т�^r����j�p<(�MX��͐��B��H�ͫ�Tlk%,Π}�y�9�b�/���R`0��a����xA���E�`�vU=�b���U�Jl9n9U*�Lѽd3���z���θ�Z�_�5��$*��_�sA5ʴH>B�m�ByP��vo_�&C~��&�W�3�~Y��z���D���%�W�Rb�^`��I�1�e�Aթ����H@�В��;\��"XSF~�k�[�^��ۙ��])h�G��"!�f
r�r��=�@��ЈQ�y�!�}K�ـ�$0T{Q7��h���� �uV3çLԮ�s�XlxVHYEB    fa00    1b30-IIpN����"���N�Z�iA
=�>�o�Y����o�Á�L�&�%$�����Ÿ����u���u!h��ͥ�t���yӝX=Y�A����[ie�1ӿ��"�Bq� �� Ks�0������<$�~ݢ}���(~
0n:W�7&k�w��Bb��B���cN��lI�[-�7̀�ZIv9]KP��vUsk�Ϝ��+�~����eO( ;��N!B��`Z�*ݮ���V��ꡕ����J�bg�y��kX\5y�ܟ�14U�z��`��,��D'�%�b袰8vi��4� �`2�&S��(��wRнL��39G_\9]H��D���}�tzGxI4&lhҨ ]n
	F3�.!&Y1��
������u��r�?����Lb��K����6�$���2��B���͹�e���4$#U�/�����Ѣ��ڙ�ά\j��E���|��DNqķa}�^�s�:�m50�0����
ʝ�z 29�d�T������3�C��BG�Μ ,LZi<�is�7�H�Q������i�m�%ً�kM��"el�A󷞰�矘Go։\��!�v
%�-I8!�@���r���z����t�ڬ9�sw'����y
�˄�c����T��-X�[�����@��U<���R���(v|�lRG�l�4:)���၊�]uu���/R(+X�z�Z�؋��� �Ν�AU�Ƕ̙��oDC��&F�����3'�ϔzKD�M�|�L�͵<~:�]d����2�sv,_��ILO��'hq����y��h҃
e�d(��iNf�}T�쓋���A$x��EyS����_��{� �M ��_��/~.�8�GI�� �ץ ~w]V�5E��x 7��X��n��J�W��q1�p�����)���i�p.W�D��{��K�G_M��Q����݃60����%+�{�0���bJQ�j��������}���z��(h�% ���c^/�Y`x��c�l�ޱ��1`�ߴ�>�K֗!�=���d���L�
���qY�Q�k������+u���ݾ�YM/��	#Jv��;�V���;�_7��+��b��������P�]���SI��TbNR�s��,w [��?�����~� �"C ]��l>�۩��S�3���Q�j����|	��L��h��`�j�B�����:��4yb��]*n}Y>�{��o�=w5�\�'{p�v���5���^�.���A���mۇ��.O~jܫ��%§F%0Xˬ���e�n#e5��6�X�8�S�pP���We p^�~Gw �+�E���o}��N���v�J�v��lM4�t*�Y �����(&�00�Q <�L3��e��+��(d�-�wp�dp���,��j�N�!�J�sת�Bfq��k]z�/(��O6�QwU��4nt�݉AwT���4��Ӡ����J�:��b�z=ތ��4m�����=�JA�ڳ�������l`U(�V&����޷����;oY�q�eN;��������`���Y�� v���d�c֎٫STe�0z}ꄃ���=׋z�Ow?���s�皱pPN�w8���Ѝ����J���F_���=���������n$g���A4�Z&P6�Fv�����+\��d���@���R��T�k ���A�d��R�1ɡh�o6\��>n�T^��Uޙ��7��@ѩnPFw+�x�p���ӟ^����M4-�%Nl��ta�
�dr�V`V+;�yT0Ƥo@���s�x�B��G�R{io�`��Vh��A�8���qV!s�G��(Wn�x�k\���gr
�8j�ԍ����ԡ�[��@�Vjԃ��BA8Ji����bDA��X�Y5�s�dp��]6����+���[�mI�>�3*uO����T ��G0DAi��6����cު�m��m5n��)r*յ����w-��RpL�^���c�*��A�b}��U��(0x��g�3��W�AV�K��IPNs6Z�5�(��f�_D>*HD�B�G�� �/��F���Cm���L*5���(�wA!16���d�dV���=>tmy$́�2���
���c�F���d��DPK�XXg+�8���������-V5�;��w�A|K����&���/��� HrG�(Ϊ'`;$�7��H��\#qG̩��I����l�K�iC����m �;���\H@��떸0V���s)�Y|P���l@���������%�^��|`��6k9�� 'u3�h�%UU���h_�4V ��T_�K>0���e�ki8C��׿R���:'���R�|e*Y>�;���X�/. �6�<���F�_�N���`����k�Q�j�c�p��������ԇ�k��C+ÿJ{@��v��EO��q]C���
�L���#~bN;PPj>1������S.�dF�
�Ix�jf9����XeF)<����ٽ�kG���T�*�`Aȳ�rX�}̯J~����U�7��"c�|��߼���&�S�1�1���и��T��E��y�����X]ͮ�Ől�� ��O���{���[\e�,t�ݎ��$n�*� ��$�A��Ư��7Ruln��5:�7g�:���7���.j�T���2��-H���6a�x|���j]mF�ž�{���]k��.�)����q�;�%�g@���%�(�g�A���m�CyB�Rh�T���m�&�z�Ě�g�Lq������:�?�ᶐ\q��Γ8<ၐYwT>�\���M	e��5���T7BJ�*ˊ�(&�u��v���9̓=q A=�@Y���og}�I
զ�!D��sN�������L��ty�'���U쿑�y����+c� ��� #cԐ���#!ؖ{���~�(n�%'�`�ӯ���9�$��Zy�L��(=�����F����.8��[�H"j\��LdYz`��yh��bX6JvMM��H�4��J��i�(s(D���wT�3&�a�q����{"T�
N����q������Qp��K6lj?q!�YRO`��,��~&L�-3t'��#�?��5��r�h��J`�'_Vp�H��P��Tq���ǆ]�$��R'�$�J��k>nL�N4����TV��>�+��wA�w׊4p`=��J5�,�Q�j�Y��|�ۊp�)��%��
{Er�t6x��Q�&6�����������_�f�G��7��r��IY_@�,�w� {��`�Ł� ��S�%M]��!ɪ�c
��_\���ݵ�Nͫ�=�\�1m�RHwA-;M�o���x���#d˪
Z��i�o	�1�r�Z^�c��[����@9c`�90���b�̏��v��Z�3���$ҌF��@G2j�)�D�e�'Q�x��Q��K� 'NO��Z�ՠ�=������&�Btf�Sl�6饽7�|�ԫ�$�X���C.M��wY��ޒ ŵ�A�O�Q��}��L�/�pn�t��������6Mw����T/ӳ
Q`��Z�ˣ�\э��,��\��f�e�ʩ�y���o����&�Z�}A��D�B�U��i � �V�U}g`LA�ժNae7����M8]㩴�RR�94��F�a��S��m'�_�;4ܼ-�j��6)��aJ~�\��|�(�����i�T+����D ��j}����SF6�/��	-�T�J�����H$ӽaySq�a���[�O���X�KHN���� �;�G��(q��՞hP���,����o.�bD)۳h�KxXMj��4	Mn�7�0=�\������ovhp8�'B��)X���xk��"%XT�	@�dD�˫D�������4��l��|G��(8MN�6�^!u���S��^�liOw =�b�0�&�|����X�i�}I}@��d��j6����i���vz/��0����Wom庎�(�5��՟�����*���D��1�`� ��G$`=�E�3��*+�=X�Y�\�1��^�yݷ�s�*��آ�����#lύ��U/^JgFlkN���C�C�S��|�Ah����4����bMe��Ѥ�A�N�J�G��NS�8(D���D��o22��r�5߭ʊ��b*b���B���rG�{��֬���,>����e��j���9E��R��Qebz�W{�����N'���x�F�k���z��M����#�C��	���%mL��9$wa�kc����팬@�,��x��a�wQ�w��*�X�er��9�n��X��jG�-X����DB�ʹ��G�_���-o�qmU��̆ʠEyu�X�8!�TYv*9���%a��� �f��xI�0�Ŗ��G 䫖��ȉ!m��mڒ�Sr�2&�W~�l�m��Ű����B�Z�Db-�$V̭�5�*r ��>�عO|oWm�����\?J�=�7{��Е���P]�(�	��gO�W$\��ea��2�FC�|��E�K�
�2�꧖�3nТ�F��n�����3�C��Id+�d��b6d���^\g�#�����5��0D`xg�y�k���K�/l����C��%L�I۾*`�����>s��G&^i�ؚB�-+"�wɆc����IKkΔ�� �S�l8x��Y�hF1�����c0~3=���X#��~1&�_�[У�_��$�<���Jty4���T��-ӎ�v@�n�J��
��HS��n�i��1� ��u�P���>���79��+��{]�0rV�t���츐}Ġ/U���<�㋞�|.ě��m��:K�3 <�]X�]��֓3�>huy��K��X3e��_��[4�#Ǻo��3�KR!�SΣy�PJ��n0���(`C)�i�O�y.ʊ�y��%v��o��M}un�s�loS�Á1ݒD:V�8��ƹ� ���*��y��i���w�+���B�@�ʵ��Jʒ�x�Lv��/�!u�,�� m�x��O~s#�X�ٗ2��_��-�;&�2������� �������<���q��1p�&y�J�U�&pց�G+H�*D��tu��+I� �D��N�8uW�"����7z��B2�c�Bh;t��v��]/�q �W6/p1Te��g��al*���h�M����SW�O�\Q����AR���}�k�b�/�!E�� ))�+2�B�9�`��e�Gȃ.�xEW��-Z��z��f�y@]�u�d
��|��j�E3bڝj��Z��j��*�����e%�Wmal�a�~���9��X��8��bS͐�;��� A� _��ձ�q�61<�����½I��qd��[|,ǘ��6�*1�@��`b$*�!�+7s�r�}MI5x���+�qz.EMi�:���W�Mӫ��D�(�QZ����j�A�Xɑ_sB�UЦ5d��)0�e�`��[K\�7w]g�1�P�f��<G���#*�c�0*N$�*+<"�3j"�z=:6>]\{��w䬉˿x���c.D�xp��($"��壬c]9z�7�]���#�y-�^}��5l��BV�G���H�i0�|�}�𜖳��,��7�J�!{��a�{��8'%��������y�%�e5�K�*A�VE!�����t��i"��zWL2�4������yW*��F��o;��f��R�XY�Ғd&����	�.+q�p�9Y�.N��x{O(�QX�58oIȺ?J�Kga�{�u��XU��q��o:8���#��K��^�83�3�%b��V���ħ���O�Z��u�Q��b(��:[��'(A	���a;�����t�4�g�q�� J�	�~���7xMPp�?��-�;�����1�军s]�!���g\A{m�U��&e{�	4I�����d�\i���Yh���l�	��NQ�#���!]'#̬���0�O����
�(+gZv�tt����@�9��
$7Ӄ��e�G$��Q�1n5U�_]ʞ�cfx�FM� �oS�S����H;)��|�Y6ԋ~�G$�Ϭ���(ϵML~���x����m[�M�]���A@�C��Fo�/�����Om�����g�`j?��
pA0N^B\�`LWڥ|�4g��Ww����UX�������e�����K�^FW[����^{O^� 7���r�)6�ۧ������U��I��+��K�]nv7'�Z��osC:����<]G�õ�ltj��ۮ>|�����I]��os�����y��($'t�D/����	�b���)s§�9,8��i����l_94��n"J��]�gh*l5u���:twLF��	ܟ�ލ]���ze�̤�� ��f�Vd��^�������7���~��cSƸ	4��u.B��~����ꗃ�/i�jK�X��O�����!��E\?�IRĤ��'ļ�H�7���d�s�u����螡!���q�	���������	i6���Sd�$z�����d�e:b�;5�!<݋5�s'	p��F��y�#v|���j��������e�ﻛ��\��L�ÒƁ�u�=:��0�"�#��� �3����1�C'kU��j������pJ?��*��'����K:݈@mt��7���%z2;�U^d���b��h&o���҂tDY[No'�SG�:�\k��%��yH�p�i�yTy����pM]�wf�u5���X�+��@:��T��@ݐE<�7�j5@���̕W�le�{
�Lv%��߫�g T��c��)<��|�����\Q��J����niܮ�|�iJ�	�ɩ��
��_@�c,<���(�7[��S3�lnn�|S׫-㎴&%C�=�
����_�tЁ�K�����7~���. ��B���~e�B=X�!t0+�-d`�5�)A��,�*��R��]ɢn�fjK,O��PXlxVHYEB    fa00    1950��T*�e���o!:$3���7�����qF�A�ެj�0�
2�k�*�ӓ$w-��}���ىq�m��PEVGi�e���f�U���%)2��K���;�y�������=�q*�(�+/��{��	�,f'�@�͌Sc���¥�~�G�y��CWZީ�{����ȥ��C���O[ݕ$Op��Ae��N�h�V���w��G���b�vpa�j�������Nw��y��4b�=ޯ�P,�}�)\��C��j�j�@k���tP�M{��2�Fn�mb���������C��9���?9�2(����@��D��w��˦Qc��k`����	�p�Qq�����
�د�>�E�]6C_}���>U �b�������#������	:�]�Ky��� �l{���/�]�-ԑ�+�Ã�ɶb2��m��;G���v���3q�z|y���s�:���N���X68��6^M��%���*Vwj=U:�f�Ǆ=$��4N��<���E�}Z5�����O#�O��mE�����vw����982����i�9�����������4�ҏd�b�POOa�Ax1�Q��zp��S�s``�qi�~��u���%�8��f�J	o���ۛ8]#�d�5d��_��r;��v�ΪU�_��94�6�͕���_˛��R�����w���7� 3]� ��st1�ʶG��\/����q��枖F�8�J�^��T϶7Gm��h����@�:sam[��l��e��R;� {�5��;�ڥ���h�|�zx�7�K@�r4��	�@���)cu�J���*HCƢR��Z�����#*��޺���&lEiL-*�4������m� ��=��ͣ!ghj��/ه��QC�h��GU��`�_�\��|f*�]�~��@�~ӛ��[���Y �N3��(���z#R��) �E��жE��k=ŪEO��yV�'�z�Z���!,.���L)LZ�<�A.�z��=̤9��\��n���駀��>k���q5KsFs舔�k���XT�H�4[����۸3�&bT�1��u\!�����0?+��"�%��w�3� ��
�6Z�8�C�j�l(�3�`�S?{� �D��W�+��Lu#Bj(3f����C��eݕ^���(>��.��7ԯ��Y[W��W�u׀'�Ф����޴�p�xa,��3{%�o�?v,j�W��U�䅁2�&v�J��������M�	�o��9��k [����Y�Kz)���i�^q��RC,R���?����5.u랚�>oZ�e4�x��v�|�hxd��=��( �p1��"��;8͇bg+F�J��*����́`\�����#�װqz�8X���%+vC���M}���g:�WA7����{�M�V��Cгe!�Br��Jh֤5��s�?g=��Q�:~X��$'V�mXz��~�Q(e�o�XQ�$+�pWW��Yh#b�����D~�xު?�Kґ��𧍆�Co�R	|�_���;WW1�ڴЪ|�N�(@��!��%���F��B�!2�"f��JB �~'����~�A��.��8Л1�R���|��@ڛHB�m�Z�SJ��3d���)�5Ď�O����-��/���I�!l�U͎v����9�΅�����|�����V:�&F&�m!:�����ҙ���^�Π�N�3�����g�sR��׋湟��An'Β��^t�����T�W��n&�0�}S}\�+%(**��B����w���&�ܬ��O��xx_��:����S2�Я�阥�����Z�XFmuZ>X��w
�oӒ�ѣ�f�)(I�ٶ�,\cvW����E�IU�|N�L��Pk)�_e?���
Y�&���-�x�g�.�m޺\9*� �k(����w����۽׊�
�WCe���ͣ%���	���pL޶ٷ�|���������%U�t��-���lcv�l��n�Ӓ�z�������3��T�7�2�U?��,��e�괊}G!�c��6m:��o|��%zZ��_O��8g]���P�s=`;kO�oߟg����cߑ+.�rw�V�`�G<>k)O=�ܣ��.�B����.�����yd�lQ��a�^�n��������u� �sԐ{�RY>շ�')}$�����C0�:����ٿ�צ�s5k�� ��KO�i�vݮI��8��jol�ҠL�<�u&
����a�.��@���?�&d����_ZQ��g$f{W�������>@G�9��p7���4�2�h� �D��[b�cK�������5�Iv���~�B�"�M�F�g���G�yY���!E\�-����� /<K�ɖW�ul�h�����sI�.E��I '�T�ҳt)�=]̙n�U�*����̿���`���4UѤ�MԂ�	�X�?���К�ic�K���s�!s��wQ���%M��e	�2I�GrgYO�HO�R�u�hqg�|���+-��N�#�)�HL�X�z��`o�]ȋ�1/����"��fK�r%c[~z�a���zr]��gZ��U�xE�ʫ��R��x�l�N���۳7yzx�x�Њ6���]8_�Q~�bL�+�W�pX
��13IP.M _/)�:�_��/Qk����zEx$��"� ��;6�ό�` #�����5�w�r��|�j,�u���ҥS`�����W����d!Ώ� A��íض�QQe�O�&8�v2R��q���r�I�����<V �>��*o;�t�֣ uy|�	��7RR���:�lB;�~	;K��lkJ��_��y���k�#7�m�/>�2��GڮǼ;8�! )n����;�7_f�j���u��M�K�qq+���y�fu�	cL�Z�r/>0vNC��J�����XrV��d�J�=�5����?ԧ����e�)=Ir�X�G-�M��ǻؓ-�5�3�#̿�����	����c"V]�KN5	Yp�\<t���i�*#3W0W�Ui�xK8���^���.�MA�A��>P��"XH`͜x5|ۢ���j�,Xf�ܝK�rWA4*u2b�5��4�˙V��˻5��A���/\>�r�9�`�αǺy��W���8L
�J4�=P�"�(TZ`%_^�G��^�
��c�-�9�C��B��_��i�ew��z�p[7�B�@�-���T�^s�t�כ"���'�����8,C���`��[�o��>s`�LS-*���+)�u��*�U�x���f�d�L�ï�BH\�s�qc��J��2��嘥����6�4�Zt�1�>R5�^��g��;�� T9�8ϫ�ջ�:�;��Xi_��r
�ԭ�w"�Q~�-~�*��m�c"��A�����S��-����	���N�O���m�ɥh�&�������oP���FYB��]R����G�����o��~Y�21����PsUo��p8qa�V���IZ�x_
u�*m,8����&�BfN��>��LGY��̶���w_u4Q�yo)gK5DQ��\����|"~���?���dBu­�YJv���7� [��X��t��W15}��M;��I.ӳ4��0�]_5H	������G��#�񱸏�����CIw�j�\��7��"ؗ��V&�4�.����
o�Ix �s�t,M�@�~��4��|>E�w�[[m��Ǩ��\t��r�6���^�6�l�z���ͮ���@��c ��S��䚏+��+vFE4�H&�bI"�W�$Ď%��P������o*�ֳ��rXV2\&�k��)�L��u�b�Z��r�z��q�J���Sn���eR$^Q>wz^��DS���v�h/��:�h��g��
�H��I�"@(�o����_���Z� ��(ζa+ipw�[�$����ޮ�Q�X��Cv�l�#��U����Q�K��˹5!�~�K��U��֤��i��e�h�fD1ʚj��R�lCX��;���8���&5n]v�ܪ�O�X�cҞ��1���˓�D͵����5�^Y��O��1a�������\����R�q9�?�&?� � ��R��SvW�ن���7���SS$�R�F��s���=���c������l����2���1W� =������P����9�K�}������5�QN ���Ԑ�����5�l�Uw N�}����ot?#�]U�CfA�=��Ǎ���AΘ=m��n&F�z�+9�@ߖ~[��_徑g0%��v����:���I��������㊀�L�~Iry
�Y��^j?���\z�s��T3$L�6�q�&�pQ��p�i�6L�4�șӋC��>���<0��ɥ@+��ĐZd7M�̸�n5]��E7�:�SN�U/�[l�j_Z\�z���Z��H���=����7��(ezx�}M{(S݈���杓p���eG�#����b/J&E����((d5�J�	��#��ɪ�8}ℜ��`�_߮����+�Z�vc(G�LU.u�M�.P��$E��(��t-AŎk!t#����y�\Dq�����������0�ϙ�[fܶ�C�D�h�cq1�!4��������E��q��e�5/��q�*�X-�jk�:=�x� ���v�b%�:=m����\ǵ���~ � I������ �jt�.�wR�pY�0��1�e��#gԖ��ˍUX��Ii6��A�QT��Lx/Q���<��R��Q�ZUy{��W�y+�\��c�$�{���F*ߛټ����Eag<l#�~Y����a	 *F����C"�
A�eq�P�8�^�Î.Il<ͱ��|5%��ʠ_	��+z��U�lџ
�P̕���;�s�����q��~��j�?]l�s��I����rTbo�1dNk8jVw�Π��C�pE�%�|_�~O�[���������Y�3k�݃�z��^TB��'�hUi���Z}��'{D�G������_I��k"��RĤr笉��4)i�04��Գ��)얓Y��~衡:��K����~��������σ6�Z���!.�����l)*� ���Y���o�Zw�	��3��~��9Z����0�E��A��wq��Ƙ"ޓA�	�1RX�?��ѽ������Ȋ1U����#���B�&����PG���+���S�5�����*���F|���	�����L�YM��P ��V��lH�Ȁ�m����Kq�~"��/��֟���^�������{B/�����Gt��"V�3c4�X��*>m6b����K����_�wgQ��1'}^�%�*U�1��AT(�6���q�O�22�^�yR�)y�{������9H�8�N��d]�q����`��2�x翱�dU����L"��?0��,�a��m��5���g�Z3�^��<��ʰ�K��e������|���4'<ꂣU1Ca:`�2P���$8d܌��% ��4�n�W�-:�Ef:���(���((��� cG@E� �@F.Z&E�k�z��{����V�W���L>��6�h��Փ":7�߰#�@eqA�t��ow֣�X%����GP���q��چ��Z+E�~z�eF��*Wof�^�s��G�Q|�x_.VE͜-6��D�^;�ӕ���F$���XȆR�Vr��<�?j��q�rM�ͳ�FÓ٩HUԱ���,���#Nt�a1��)�P��ٗ����^}�`�Y���՗<��<GHi�U�߾���������y��7��}�4�1O���=�BH�d_'��'��3,Ux�� ��M�_��(�:�J�#E�מK�}�9�w,|yu|��iv6�&D%��&���cJ9^^`O�$�G�ҵ���z�U@�T3~[���fF��ic�9��|L43�E5c�cy������V4�y�#��.��(�.��xB�� =�����\�9�T�X�|�K�|ɺ�q� �e�؀�z���y95���=�a���B��$aÂ��d��H��{��3Mn
+6R����M]&z,�}��8��>a�vK�D�lv���,m�����k
d�gX %�x��z(L���7)����r�da��.��گ�q% �a&t��_l���*����� ��P�h�%��uVϾ:���KP'%(�h9��Rkp�
��W����8H�q��E�[Z��J8��aLw,��,���'DS10v	#F�������ގ�Aq�*�/� ~u��u�-�v��;�S�\^s��X�rJf�Չ0ܓR5�����i`�e:3�1Xa�i֦Q:ZU&-��տ_mr����@u�����d
�*�x6��3�&,킎������ߨb���v���F���!��=�Aڧ-63TJaY8�~d��IPf��퍎fRE�F����
{�3�A�=5��s_�Ry�NQ�e9��XlxVHYEB    4f27     d40�&����w� Et���J�PrP�!��g���S�Y���E"p�H�R�Q��B?Q�Ȗ!=��u��W�Q2����5���v��"��ˎ�Q=�j�_GOk�(���BX\��WxbOS�{H�D�d��ۯGx��?�6n:���y^�%q�p��k�C��%���	ȡHx�=��Ӛ��6�a���k�&5E=��}�0o����U)�wX��SO;�)waΫ�Z��:=��D�~����j��C��sXj��@�\�G'Y��S�hpp%I�=�:�B����D��)x�u
(�k�\ ���fm8���a��/'T�*=y��5ė������c)�*e�����:&���7fI2:�/�;�hZ��:k:�@=�	�̪7�XT}�����f���UPz�"Z���;���t���$�0V�\3������#@�">$����!����Q$׈TN6�0��a�=� )?|�G�؈7ʽM�YO�>�'��It�A�@��n
�w!CK-T���RbL�[J΢�0��X8�*�1qH3��>4MTf�ޘ]���z�$G<'�r��ќ��c67c��nO%���9�R��SX��ڰxr�I۝��4KZ�4X�|�O�gm�}�\z�\Xx�"ׂ�+����Ŵf���<P��K(T��7fJ>r�:8�Rٗq�؄ps�g�*d�,F�}'����~��^8����(�eM�I�T:>�5�}�I�v@�������%_�(��*�bɶn�]`c�kdm0��D�Ȑ�"�K�גC�0��]d��O���=�tpƟ�]���]m�L��nUO0�����&����{�����7y�q�г���~#���a��5� ��*�K���8~����l4Ө�uUe3~ו���k��&z���j;����M ���?�	-�&�V�M
�s�QK�4 �v��|�5S0��9���������!p��M�1�WY:)����1�@�@����������K��lm���΅�Ѯ¹>D�&�r��m��Fs��P�\���"��H�^KfQ᜔�dA�\���@G~A��.�-ZMS���P�gF3��w���x�`�J��2<h�úA ��D��rJԸ���V`(�:�E���%�R����ؘ�&���GS���;�
k�3���$��2����	Dsj�q= ��s/#ٷû
���ow���Ԃ��^��p#i���ҙ�og�P�Iz�^���Cr�R8亦�����Žx�5q�f��&3b�R�li� )�J�7-_9w�S�i���(�V��a0V�#��/�_~H���fC�"V/�e��h�du+�#�FW6ω\FK�Ґ���Nګ�e0*�S����/�62��(�9�{9d����]-n��ϽE#����.4-lJM^����F�N���v��	[���+ͮcZ�,�N���Vt���Hi������Did̲���+[=��\�MQVĒ�����q��|��U"G�zk��V�ֲL+����r�FN(�MP�yc��!���^�����������C�h���x���/K�2��q"j '��)Y�$o���5��+>鴥OH>#]����R�!%	���4�y5���6K����I����ܛ�e#p�g����'g>̯TOLr�����LT�P��2b��'F\���ċ�'��>�G.#�$As���UZKF�N�h�Iǚ��$��ٿA�<���ۋ^��3{���0y2���z8=�����H�-�g��w/C�!�q��$�9
�n���O�6�6�qHU?�H�i�,�	�;����Ӌ�(�����c!0j1>+�.�@�[>�.ۥ��m�U�g�v����B�*Y�W{Ϡ�2�>�|rh�tX[[��d�w��)����t�I���~����t�K��ǔ����!*S����b4ӟ��=�z���N��m��Q%�a��cD�������GV[^̪�c��]A��q���p��/h��}�5�2����u�S���;�jߓ�����y�E��%�ݲ��@p�!562�o1Y�������
��J+K�F6?g���agU�{����]�-�.�N���^���D�J?�j;�W4O4|�a�|�����2*�f��ҮR8�$���Hx�g��`CC_�C�q��=�
��~ŏ�_�Yw@|)���kK�'#^��@��c����T���o��_��a�joV���b�:}S1ϫ��i3���������どZʱf�a��
�.t�}̳M��� n�K�Ǭ)v�}uJw�9A,[v��iψ��.݊!�v���U���l��fD�&�7f-�ڭ9;O��N'X�������5���A�9�>�c�����}^��@��HNZ���,'�If��m �Ɍ.�w�fE�a�T |Tj�cR߂emT�v���NL���L��-�l��A�bs��Bk�
�����C�������1�!/-Dp�Ҟ� ��S�����4���8��s
�bc�Y%.����z<���T�b�6Ö��"���֞±XR�-˦�V�L�ե��W�N����e�;��7k�z�Zq��m��X&�U���9C�Gv�[H�]���0��nc�{`���,e-����y�����]�u*�|(�M�Eѭ��dQ�j��u��s��E�9K^� w$�r`c���˼�6V)�`x�i����%ljb����K��h�����N��M�Ih�*���E)vS�A�%�3���+�_��$f���ky�:+e?����o#Y�o�}��u��l����{x��+2����DMA��k@��s�We��m�,1�G���o�	D|h��F�ͺ�ٯ���iSnO��ͩ?� ���G���y�,N@�}r�,\��m@����wކ�w!<����)#TA�K�����^�G-KUdU�`��Ö�|Y�sS&�f��{;r��GXׁb���`�}�aT-��]D �3/*�t?���+Cޚ��6.�p���+�sm7�aGX�0���q���E2�h�`(���»��s�^��3Q�?Ҹpw����j�b��G���Z�a���|��Fɏ6�+��)vѨ���T i����S�tB׭b�&�b��M�v�'�����3h��ĕ_��"]!=2�W���N�zn���>rj�`#�KO'=q�������O�Mr ����h�;�vM�]i!L'��Ъ�?1@R^�"���/š�jg��b�����k/(���R�QΔ�� C  E��/��M6k�/����I���d�$�]��1ZG3���s�OJ����3���T!�u��