XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:�L�;��Upk_��b�;�X�"���J����Ȩ��"q8
PB�[۵L�'�u�A�	�=¤?�)#����y�����d��<���~&���ք�q�-�|m�+(�H6K���]����N4.B���j���P��k}�r�>�lVnC����iE<^L����-_�yR�����C����1�g���S��l�k}ov2�0^<ᑥ����6��9]ѽTU#`�tD�+��� P�^P�+D���!�ƌcS�����[���c��c��A:Uh"7��i�к �}y(�҅�C��c�����+�'#X�C�s�#,9�/$��ף6�$v���8L��+�s��e�_��k	��sk>26��'̖��x�1�9۪�`2F&Q�z;�qy�gi{�:T
&@"QFT;=/˪-��4�q�:Jǲ_.V�G�`D��.m� ��z��iq��D��Ū1�/05y��F&���}6�0����?$p�if�R9�m%

GX@5h��\��q���Mn���H[�Ԡ��xZ�J�B!"\�K�Ri�\�3��k��g'�����0��;�;�}d~�j�]é��z�H��6�g�#�����:YX q��͖��$�����M��@v1�����Tj�QB�/�$�竊�/�+S=��T�cS�k��94��"��m�>urQ�`����īʱ�I��K�/���OƤ�c����u��3ن��@j�;�.��n����t[4a�B�;��0Da?�z�J���XlxVHYEB    aa52    13d0<��[P��v~ii h��s�8|d�\r;�q
��K��4��3����P��/��&y4�Ͱ�)�P�$�L0�)�`쥵\�{ظ�66w^O��:>��(rS�>�=���k��g�EE.��D	ث���k؍��jJ�&x(���QP���6݉N�Ԗ
W���*>���Aa���\,Nc��v�v0@o��>��6��n� �Ҏa۶x���kė�Ł���g�!�NlJ��uM~	����V��RN��+��7�_Yk�C�Tk ��J$
>��߉<���l���
��W��Ńm�͈r�S�%\8?���B��b�[�:lE���4��#����� C�|	W�?���q�W*���w1������^`�q�F�쬖BX��=�%b��Z�샂F(���dl^��|V��7{��D���^�X	:!�G��?Ѕ����*��Oz��L���u>d��3nߗ2'0W�>���u+Jȑ�r�Gb���;���[��E�[��P�Y�����p[ԍN�BL�L�G��������]�?�£�*�ƕ+�bh���J	�sO�sY��ay>��)OR�:!p	7b���h�jwW��d�)	�}� ֎�Ai.�M�]L�VW�;�X�77B0��'\@8'�:��ͳd�u�b���}��@�O �<^�,�U��2��'�����@U&���2a�����p�4���0���E�#n�c��0jm7h�:���T�c�����=���ִ�oUe��o���D���:r��I�3+o��Q�.����.�#��u�)|}:g)�E�7>�kެZZ_��*Jδ��4���B��I���T�0#�#4hla`1�2̻h窭�F.s��$�d�JG��2�0�5�����4���^�?�	)�bT/�%H'+�XP��J�"����Q���ap�~��=�~M��w��?���ʑ�K0iTb}�^�Q@JX8c_2Z4A�_,h���cd�����7e{���S̛QꞚ֎�[ e0R���:ne�\[�����!���c�L����5:m3X�Q�k�9���Y�1�L��'�4l*ue���>��w���#P2;�h��tr�J4���Y����5Q��m ���\�s~�
��Ix���de-�k��h��R�v�U�7�+�K�NJ��8��4�%u�)@|#�_p��o���  ��|���E/�S���<�.E<r�.`�9^=G6ڽ�RD�@�to4���-���)���W�;tdRw�<����)�|=Q����@�FJxB�$$%�&_�I�u�z��Ժ����ivz#�I�y$1�	�c�֤ú�/�h�P;���kk�_�����w܃�v�o�֡ImR��}D�$�{@u�!��:�o�B�)�H|�tG�$y��;�sc8�X�!���"���L���3',�J��(��԰h�<�E�'�(�~����.lD>� 1��b�}�y�Y�и��!YO��.��Rٔ��d���;�0-1�Zr�iJ!F!MC�Z%}��2��aBy���Z-U�yk�����3��.;����|�[<KמIotC�+��?�D^�	���I�3,'���-|��1�k�$�ɤ�L��{��Z`pC��z �^�t��=:Qu�|�"a%j�;������E��ܿ�K�����dyT7}E&]��jf>��n�jR�ܬ`{�`1�����~���eX�����E��� '�:�m��L�k7�H��/��9��*�}�@�)R�f'R���0/!�K�8Z��67�xA��wS0�c�(�@#�׏RDK{������@�z��%��Kl�q���0����#���]�<E�f���ǩ6��3��L &e6xj5��9���^8���~j�$�V���bW��F��W�����g�dś�~
G���k�I�7��f�F��E'B�|p�bЮK��"�D����v�"�y59�.lQ��쾲�i`��u�`������u[M�"��,3?�'pՄ��E^�z-��LH`�{V}�O.��a.ʯ����{t�zN�2�ݭ�gѹP��?J���o�0�c�8��ʱe�z�sj}����VQ�P�3G�>�&J�B���/9��.�
��%�~���3�5>�n�_9�k�p��}�D�/s8 Q�(���y�?��Ed��`7��=�@$чM}ɏٱ\A��eC�l�=(�b��B(���I^��x�����پ f׋��
%��X�1�m�mA�M�w�t�l�N�e,(z����+S�iFA��E�=<Yi���E�S���,�Cw^:�ȡ�3��6L9�R�͛(ۻDu�}�E�� �Ѽqce�W���(�8�5��;�`�r�UA/B�2��eӒ}6�5q�9�)7��>��:v�C9C��J�s�7���,�3�OF������!?�i �8Xu0�7��d�wR\y�⍇}I�֡������h�+d��c�b�.�������$) f�, �ٰ\���,p���@��)gy��E۠A��bQ�
r2�&t�[�#��?���w{�B4	2�M�}v�O!]ȋ�_D�%��V��l��6��A4�_?�+U�$�s:9�j�Y�"1�ö����2��&�:d���C� LQC�Q�zB��|q�r�u����S��O�"򆼍�n!ɂ��1��bh����v�{~h)ϴ�=>g菀xP��u��Yj\*�o?���=��2w{澘y%��Nw�N����t$��ɖ�{9����.
�:;�)��O۳8'�q�f=n�����∣=�8ߊ�
oV
lDc�2#�Q'1]����`�ħ�q�-	n$����]޼dS�2�R{��֍�o�ofk�~�v�Ռ���Z5/�Q%����=,�P^m]ƧM�^M��eT�w̑��)H�9��@'��C/��'Ս���Sjok���U��1b?O�ߞ�@E�ɟ�?�
��t��<Zn2���D���&M�7����>u���Ϛ�L�/V�p�X���?�lx���V~�]ē�HnAY��+�& }jS��j��g�:����rJY*��;��E#~F�
��yOHc�Nm6��� ��{4(�
l6l�ˑM��1X�WҺ�*eUy\�}M}x*@݄�9��΅#N�z�	�+�!=�]���0f��͜�]]n�ޢRh�5S���tDD�P=����3<:g��!��� ���)���?' �sGc)��[&\�JW��b��w?5��6��e��Jg��w������S�s�k� �-�_R���HF킍Ψ�０�'�&����З��0K�R{����	�Vq���i!0���d�Q�@ʵq)'sB@�+nS����'��'��v�7���9K�����������L����0���4�1M��,���W����y�L<�I¶"���犎��kҡ0읗R�)n@�4g���Xr.�A�+�u�Xp�i1�/sC�P�i��*yX1V�e`�׻�r���6^�F�
��HC�8HTMHEՂ�J��) {��Rˠ(3����P�"ñ��GA�0����δ�kp����p���]'�\���aj���%�(�`��Z]�=3����ғ�P���u��Ŗ&*��u��_ {<hFV"�p��<p5(V��>R���|q#H�S�>�ӊ#�矕�ƒ�<��ʙM�Y������"C$B�B���8�Ѻ}�d6GM-|�W@Rj��d��>����6�o9F%m��|��iH�MMM@�T���DԵ0<���>�R�l�`�A"�{�B3�3��z�_Ac��kƈ�O��ht+�ꈀS`�.;[�T@-� BC��Tĵ� �Ux�p ��v��[��C%�a�M�ӗ� e�p��������'�]^�]J����e�Ϋ0� \���ϫ\eLv|���B�ru��-��DB�����y=a�@��g�{�Ȯ���-5	h1M2n8����谯��;3ľ���#�Z'!�&
�B*S���`����f��Ʒ�-C3�}6�k�*e��R��{��YC@<I�c��-[�M#���R=!�I*��U%RŢn��֝^NT������p���LH����B�8�!Q%�O35�#��T(Y�F����2J�����G���d"f��,*�`Q��*�ZC&Ϙ'ɻ(�s>�iӶ4�@�t�����g���h:�!��%���[Sz�7�c���8�!R!^������W�G9��}�#����`Y_�EdyVȸf�'��Iq��2���>x4���}���y�ȧZƽU�u�)0��J���(��`�q���E��'d��wA�ĈͽS0Vs4Ot2�_���qPL֕h(�ğJ�6�\v��qY�S��}r#e�Ә� s���$?��J��5���h�G��Z�
zO������s�o�3p�~ǒ6����F�F�!�PɢµXք]E�S�N)����3f�����\��0����vѡY#��DMҵ9���W�Č6�h>|�l2�#��$ƺ�2Y�QU��<$���0�h�d�qyS�`�bf��n�yQ�C�U�ܶHA�*C��A�����5�:�+a.��a��PiaJ�(WEH�!��)���N�V�ib�q�#vX�bw"¹:���r� �! %ʫ�?c�����8��;*>���qͬ�F5N[��#F1����#��O���}�.a��|ӓ����d{/I	���ǅ���L�B|ܼB*��ݓ<|0t����-Ң�|�k�}���#� �|L̀V����n�q���G������Mw�Hٸ]ܡ���/p�h'� H'���_w���7�J��E�UJ�I0%���5#'^� #I#�i>�n��O�]R[7R�P�kC�;��$��BvR�z���9�+t?&���7�g��z�8��^|���]��rHfR�i�c��~��t� h��``4^̆0h��mD�:-��3�I�I�<8~�p*�R���š��	�����_�����	����'\��o��L>�n8��z��V�3���V