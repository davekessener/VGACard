XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����`�5e��93D˲A�V������d#��Lb0�Gˢ�ʖ��ۺ� �����Pc�Me�'ι�׿�|��O���T��\(�t�H}&����+S�
�0�ȁ'蕸B�����Q:���b�q�����\O��:rO3�	�ʆ��K�C3`���<t�j�F�V���i�3-���&��P*bt_�?���D��j���<-�p�����|�����\�3�>9�3����l�sp9K��,K�pu�U<�uA��j�s��3A��fB�5����Qri�#�-k���z�u�7+�ؓ��R���Ѝ��!kTn=L����J0�f�BWD����UӸ.R����{�9B_Ӂ��?5�(1%�Z|[�8�Κ?��"o��_~�qJ�mtö�%���M��ʪ�7��VJ+�����s���N�3�Mx��3�'KR�����'ɳ��4x�b�'Ґ0�1]��k���Z���j!6��݂z_pI���H�Jk@�y�����6[��ʠ��s�'�2��b�>ɥm�d�ZN��)��A�g`o���F�֌���L@�a�_���B�n|ךxfG�����SÖ2m�K �����xv�}mN�D��$�j���AL���H�ߐ!�r� �Zp��*�O�]�{������5۠� p�+|��vM��Η�/#�I�>��AUΕ����� �8��t}��3Dr�$��M���mm�e_�J`�#����mp�sc�ۇ9v��('�9�	�$��P��F��ɣXlxVHYEB    aa31    1e40�����e�
�wt�x�(2�G#'	R���?�h|�c�eŠv��}3���)6E9Ƃ��h��f ��(��`�"�S��UZ#h0Y��3E�C�X�6�E5e�S�FY�f�I�TY ��ϗJ�7�wH�X��E�yHL�
_J�vR�p�58Y�2���u�x�����|<��#�!�"�Y���b�8=\�����Y+�	a��׸�^E߸?��0�6ӺdS��m�Cρ�O[�2�: i��MMۇ���.����a��N�G���ē�W��3V�}�4�ڨ��t��E�B:�,۸I�.�����xv_�u%@�[���a��X�4tpV�we�}v+X����
���@� ݦN� >�����Υ��ٯ<Pf!�����?S>��2�׷d�/�"A9�d���.�bR�f�K�V6( �r����A��`?N��{~(WXo�׉�"�	��_�M.�o�[6Z-���dB�e�>w�z)F&B�) ��H�u���Qƙ�Z���Mx�"�*yZt� �Z|�ѭ��ˊ=9�y��\L�dB�ϴ#ы�Co�Q�ܑ��1�S)�� "n���spiT����"M^���Z*���W�v>�fR��X��P����~���~��ᰟÆ�}��NR�Yu�;H���x)�?���a&��@�tX�r�3Ȫ���A8�E�Uu9��G�N�]���p�r�_��Zڴ��J�	��/ic����B��-l��;F!�418Gh���d�����f�A��JX��%�tb����BG��5B��9"̟��s㚯o˷���B�e`/��;�a ʰ��+p�eW'��'r� W��.j�?_�6���"�o�ļ�\Q�3%:<,<T�r���%:�8�P��11|<)��d��fs��vnm�E�����K0�l�1yofq�f���VX�.r z|dSFP�n�R����]�os�������Fj�Q�f������*��)��{,l`�Y�($L��e�uX��*I�dV5gP�8�DI4ډ��Ԗ����$�P(�w�L�ff�rh`�F�!򰮁mj�oU�tt�`.�?߀y�p�/�w�9܀i�36rN�Ϙ$AJ;P^��z_Ж� _z)�j>td~�L��^�YCk՜�X'�!��1�'D)3�����~���2o���YEꥩ�f��T�7*hhW���H�e�YĜ�&�|X ��bП�*�Q��5L�zyT  nQܷ��Rm�ϝ��

ɴ��x��Y���wQ��b�/��
��LF\)�d0�hY ��_	��rc��+�l��a뇧���f@E���9P�eSJW�z�C�A��{�$z���>�J�!ݮ������Gm���*�ت+�v�Hso⤕�޽ƜT��̅e�jn�VsPN������=U�9f�vb��~D�x��Lb�Z��`�bͨ���$�DԶ[Lqw���>G���@8�Jhܴ]%�3�`��R$�c8@uY0b�5N܌�����uJ=-�DŚ�n��N��qp]x�	�c��&3�k��̑E�o�b�x��������b��<��
+�/_�ϋ�vrÛ�6�c���Q�Sb7m�F7|����ň�'���[����;[rw�P�i���<�*�����3Z���d���������1�D|�@�cU����TO=���6Ůֹm|oH�]�Φ�Q$��DC�+��=-��e]�;��-(�ۤ�S�X�7t�����c��<���󞰴�;��O��ٵ��T�Y��m7��I�$hUSxJ�q���$���u�p T��Fj��O]�
S��9�?���GM�U)��.�>8�|�|��^X������b���#�a��o)jI-(6��]�.��A�c0�� .^����V}Ծ��ˮ�>I������ǉĠ?/��`2�jO'�_���x
~�@�mgی"�o�C-�џ+�i+ޜ�X �����.�^�]'J�$۳teҙ�;1
�h��:��JX�w<Tf�T���%[����ǳ�Vйl�d�BDGZޙ�C���	���j���^�7A!��㜴1�4
O�Zŵ�1��T��H��۽�2+^�d:\�}�/"�{�%�	�>u����h#*b{c}g�����#b#�IZ�����y�[��M��a�XS���餽���3�:#�R�J�`08^�>���ԺD�S�i�j˨�F��迁��v�5�:�S7~�q��-<f35�?
y����G��R/���<�o��F�VL�N��n�3��>�[DZ[c}u�4' ��RA��`���t� �G���\*�U��b#���;�ng��mt{��d���Bs� @|"~�s�K��j��B^/ѿ�����U��~_�*���o�w����.��RS����q!�	b�cz�Gf����,�S���v=�6���7q3�-32�mU�W�4:И���I4������jܑ�L�\T���ls#���ǻ�[���c�\��~MI��kb�b$�@U�=�N�S�)z���E��/��V�Ba�7�PF#��r���!��"4�z�����N�u�	IV���S5Άϧi���DT������C?2�?�s.� g���캹��>��b�D����Zyj�V�h(ׄ��<�vr��� N����������|�\�1�k�o�8ןDU�� v#x��L��5��~�Pޚ"ӎ�������Օ *��Aq���f��+ZPi��g%�����%��β�.~��[Ħ��dB�U�m{���vu��w	�xbc���`��Hh]v밡��������Wzy/@ �g�7�s?=� �*������W?��K��Ҝ���/��W���q0m�Ȭh��l�ٳi��z5lg���$yO���e��@���)Y�s�z�~�Y�?:�������AբM��8�ݝŏ�`S�n���'D�%}([��!�� aôRP?D@_�3,�J�oǵ�`�b9����1���D[�X�<	�I]	�4 �
�����iS}�p��ѱ�^T+gt���?�yz_��#��/����A�7U��||���+Dr����z�F�]��CA�27Z]@ �� ���Թ/�ҽ���q��!١��*�Y�&�J�u[@I^����g��䓪k�S[q�c�`�ZV��=������Qr͟Ǌ�Vۈ2�
��tGͅ1�B�(`8D�5کQ�f�O6ߴ�ݓ�o����\ܷ)o��IX�%����:�JQ��ec6�����dk�1�-����l��<�ȁj@O�(��D�Nl�JK�O9וz! 5�L�#�|�s�'��ìU~�^7~ŒU[�?�ހ+7"��D8�r	��,�k�a�DقδZ,����}��o�O��t{�����5�wy����E'<����w���~����9=Z �;��LI0̐������P��0��;5��]i;s�;��d�_�j1��k���)7�;VR�=����C��O`�Lj�Is�+#�����ЀJ�������^f8�j:5W�\-eó����ϝ����e��Y  o�!; ���>���䠑C�nVyPb�>>$�߶�L���m��&��nf��{��e����c�c���Z�&�%��p&���|F{�\&�� }Y�.�y�D�j��}�H�}'d�r�h:�f�%�Ċ��q�;�zeQI��G�t�W=�x#��h���s���~�D��v���Ñ�I]�k�R�����{�E]�_���ԇ{v�`�B�����g:��&�����s��d�Ş���g;��	��s �H/��;֧U1�y�K��8@�-�Ǿ�g������lYR��}T��	���.M-�Q��_?,?�G���*�j"�e|�{�Sn�]h"]�词E(����/�D�F����\���b7Ev����[�@��	(�<����j!�;]��_�h�$���u�~�̮�J��`M"�WxD�J�(�K/D�Rc�i�=���n�M���n�o�l�<��}*�����m�L�.�\9�Z���ژ5����-�ʥ$V9jp.���k߻�����=F�V�} 2	dnP���(7��+bX&R^��$���)����D�?�̸��R�$�?�"��A���GŨ됯���_�V���W��� �E\$�b���4	E�B=l1�q�+��v#H�0-I/~�Q���t����FC��ɿ��iW�+%�(�$��.�f �`��̿�ιo�.��{3�x��1D��v�� �V~�%��	"~�B�d�Y�j7|ZE��j��; 5��#֖�DK� �{�]	���ky��rj\!V�{��:* ������p��ACZ�
�P\���1K�w~a�cfR�"�X��gfb^�\"=��L�r>pK����R�:|�㝖��O��n��i�K�C��!IȒ�VW���5^-�`�T��w���r���@Zv�������d��ˎ��9��=4��;`N��I�����T�n���>9g��,�ب:�S�I!�T�(��ꂠ#�x��U��G*l��H7a��E�m.e擞��$#��L _��$�K_��}�듟Ye܃r���rώ[-3)�H�Y '����]� %do޶*Wķ~�� ��/�bzBT4�u~��1Xi�;i�NZ�I����m�2��@:�������w�	G7��բU�p4�3�NQ��U����M�v���Y�Eu�̨Y�"rU�������U Kl�z��!�8������5�sS�M�qfBAf.A��'�'������
=˲�D4�HUpK5��Kǈ@M=�U�@��K 񄸗:�UqW�ޙ�w��BE��w���w��V�i=w܏)���T�)��c�>uq3�5��ì�����]f�!�_�9ވtkk�j6v�<���dX�(m��0�:�A�Wi�*6V�Q�o��=�M�oN�-�y��`����/���z��M_���rޣ&�'�Y?ĳ�� ��l��{�g� �W���e���oRf����H:N{�}�������]{.0���MIT�Vd�maY���0\�9�����
�wje��[��4���C�k�L5�=.oJ��SaLW�&c��d@UL�� T��s�Om1AGuB�=[�7{ʙr��w{���l�u���ĥ����y9Tg+�ߝ��u��r)�cn�|��ձC��g�	��][C�}n۩�tL�ĸ\��^ �X�!���DfZ�Nn7�}E�D)��(EG�!����?�6�u�)@F�
��$��f_��K W< �2,�(�;��S#�|��$A_�F.�2�M×jB�����"�0,˜���>��U����1Z>j�ƻfV�1��^��0�F��P`%u��K�J ��#�5|A����v����:����7���K![A��h4��gs��$fEL�\Үnϳ��.�hdƢ�����t3��B� �Zr�Z(e@����,�&{Ā�<�� ;��W"x�t"�(<J����,�^>�$�n5�T�X�*�7��M��~+�w5*�(���?b����'_�.��w���F��k\�RD6R-�\�������Sҵ�!��R�_�/�!��~������L�����A�|�bR��\+�=���K���E�o�((�?m|���W�T�Y�M�*;�M���'�Bl5j��ӰEdU�$�7o%�@��6�z� ��E?n�,�[�@e4-�����1����N�)�X��*�HNOu��������N�JK�@�1����Q�B�/��)�.�5 �/�����p\J�p���O��w%���1�[�:��1.�ҡ���)��ʴ`��¬�#���eB��V#��EwB�~��FU�#�v2�8�ZiJ���-C�A�xjoi��3 QO�%n7�5,��7��v��p��J���1��l��]cP+�W#KR0�p�h�v��L�$�g��H���	@CW��K�ir��a_�Cb�á:�<j����� <�=NA��^%��;7�����<$�����ۨ�	_o�w;��V��W(��?8�2��\��M��푻��ꡢ�g��k��XR�%q�/�-�nwU�{}�����صz5(�״Uл���wʘnܷ�N/ɤ?9�\π������|n_�I���<�UVG��*o3�GtM�_�}�P�01ŵ7�'�Z��b{S��Gij�8#](oKmoKS��UE':xeG9�
7���i�����3Tn���@��i��D!�.1X�m�M�XG�U]˙z�?S.�\�:�I�y�$���AJBpJr�^���P�:���7�:�~5c�����ac,�[R�'XŠq��i�d���i��|��������r�K0m�&�/3�����>�O]Ed�+�(}k��/|��*�����u�x(� �M�X=���������4�S �Zm�`mD2��c�i,I�4ë�{63��h]��,t|pN����������
�|�e:D�Z}=D�+i<����e���v.5�V��1 ��Φ�8N1�`3c��r��n���M钺h��� e����̊J�����z�i0s�$��a*6d���������D�&Br�9��(��ؿ�@��#��>����@!A�������R�H&�Ӥ�mj�����w{���:��O��_m!UdHV?������J�k4�&��3�>�b�e'��}��V~d`x41��)69���nz|��D���W��KR��1�HU;WJZ�>�+yj���I���Q,Y��A���v��&���������
��Mۏ���$��Wƾ%Dc���
�<�lϢ7ʝr�S���^x�i���[�V�y���2 ɕ��vK<�@Q�/p�%����bk��c���~�Ho�3'��u�|��%����?�����;�ve� �Gk�䕛��NИ����^�;����3��\(c�?���1�L�Z�`�*^oI 
84���Plo�[���|�}�ě�b-T���� q;I��s;��J�u5ኀ�\ؕ4�;��!-��g
�у�.@_�3��j���͎����	h�{�4�ג�:.�:��	�X*9�Ht˸��$
����o�*�L�gq�����"�]�-��������ʃ�a��Ks�( �_`)����lP*6�y�z	��';uw����z�����c\�17G)�_��b�u2��~�
ݳ�b�)���x�������\䒃�J�m�a뷩xA{tD!�x�����H� kP%��ҽٿ���i����OB��!K?j{U����9�����ɨU�D��@�4�Es�hox�B� g�7��t�Ŋq"�4F�eʞNՌ5 �o�����ј9�{��3t�B�(��h���G�-�7*���]���`u2�	��mEB
��D�W�v1x8���g������6?<��7�,�.�h�GU�;E�)؎�5$jY�t4m٪�_vB�&-���������%���!��_�b'm�秷���Fs@:K�&�Y��R�n�B�F657�N��8�Du�A������)�"KS?'�k����L'J�v��)���J5�N�ҧ���$���v ��c�L��J�����U!$iϗ�hqF�ط�ٌԴ)Ÿ�Պ������v���f*u�YS���6��