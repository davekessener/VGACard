XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���W}�N
��OKY�ƥu�w�|4�s��d��MWrO��QR_d�PT���P�\�r�[&N�2�Y�p �0�9�~c��x`�J�u*[�[��"��X�'��X��Nz�����<lc��@��I�R/	S�%�C�@_ �m(o���I�$IF�����"F�5�P�)]d��~f�U���j
xn>�$��Ʀ��#��A!&)K��4�:&BB����TPw�Z��O"�ϘS����+��j7��gi��-�:�	�9(Xz
����zc�{��O��&ȧ@�>Sv�	w���BdA@�^F�y�E�]�b�h��Թ!���$Ѕ�[dR�Ǟ^`w$��ɘ"*� �������# ��bl��f��$i{�HL��um��YG�r�kc��E&1#@��i?&��m��^�Z��:[iǓ-�a�o�nꢌ�uO]��|��S���1��ܮ�5��j=.���k%=�J�T.����B�>^�䘘�mb6J�G��`��lG�P�5�Mh�R�jO*{�4wg��
̷2
��-G��M{�vC\P�e<B��APk��~�L�Y.v�)���S�>���{�ᜮ�$�w-���r��r`�����ӓ��Zj��h-,����S��޽"��T�\���l��N&���p�ع"q���3��1y�P�e�'ߝ��g�@���wk��
�U|?I�Ե��6Â'��J'���
N�<��=�f� #��E�v)��m��S:,��[Gu~
M�b��`�yX� ���XlxVHYEB    9efe    1be00���gh���^��?[�	������5�V��*�k	ݺ�lOѮ��m��m@�*[N5%�w�g"ct;��Z
�>x4랉�Y]�^�=m�V�_{q��ӢF��D�����������OZw�21xs����	�J��<�#���~�@ݓ����/�E�9I�z���R�"Se�ݧ��)�7eʔ�W������|�a1.�q�\|�~�1@T�}��^aWb (*���}��I'��Z��� ��˰/i���Ò����Kh��0Ϡb`���e1,�Ń]�!�`���p�.�M�874�(�v�/:	��׾���a�I�h��%͝:R.74�	���%��e��\��z��JX���S���1��!U}�dj��aQt���bB�'S����hhY�<0�K��_��c�{!���'`��G�;mB�LQ�a�BA����Z\��{Y�a�$t��˿�e=������[��_� �q�&������$���2�SzE�GI'x�$j�@����_� �aD����e�^b�d�_y���\�n=��	�?oH�:WM����&�:�yO�Ԕ��h",�M�ˇ|�����y\��#@�`���L�o/zs.�<HOФو�θ��D�4{�a�6t���<��_��t���]����?ǏR�!��8͜��/�z�o�i$;���/T紗�����I�HH¸:r1�}\�h=���w"�5]��A���<�\�9��*��~~�jĢ�י���".���6��T~�>WĭH���E�B�|�����>�񪒡��ϫF�����R�}
5,�����Li�F���r��Ao�j��%ğY�|������:~�y ��X&,��i%G��l�ƎO��^GdVa0���MMo�̚?�D'���
�ě+��H(�g�І��Q�
�(C?����@���0�mOn��x4�K�v�E �f�jR覕�Km���rUG�h	QF��o�v��dbR���@+�ǜ۾� �(ĶW��h�M�����u�T��q>���]�� �w__5��h4=�Q��	�͏����z� ���`,+ݻ�1�6c����֚`��4G�GV����d�	,�T���0g��
t5�n���]B#>b�:�^(�m��SL��'3;.f7x����%�"���|&[����JV\1�I�R��Bu�!٦��q}�AK1.���bnp#�b�x�[��
>aRP�0�%��f�E6���İ���2	�t|��˛➎cP��I������{���%�Sb�Ε�
��h`w����RV� �p�7�
�bDN��[�
�
htbj��su�*�*�uqǉx����tLՏ���jtqF�-2�D+%>��FEa��8��Y�Zy,��`�&A�.�:�\�ܧX��g��Y��ɓ��6�'���/*>�Cy.�M'�>4y4������Z�¿�n�
��a��Pk��N�jI��Xv�&�K���#X�����z��憐�s#��G�]�w�E��ه�f�z-M����s�@x
#	�J�^$��*��w�1�ߦ*��~�s�.�m�ewLt�(b�L����LCԇ��h��t?�*9�Id�X�r<\����3�����������3��H�Ԣ-F;@�W����B3EH4�/�>:gWD2 D���^�n{��3�M�u52J�K�6V��sOh��4�F�x<���Lu����%�:���) ��=s1u���֘m��U �Hw����t�P�{�׳�v����hp��g�X"ot�(��P�;���!C_���f���j�]������w$+q5{�ڨ�� �ʸX�t����;nv0�)�����t�Bă�[2��מ���N��<���
�MIܹe@'�z�u 5=b�a)	1����Xe����M=
��{}�?�Xsxay{�'e��vH�te�{��>4�
kn
���&����������[6�B�!oL=�+{��'����D{<^W����VK��)�;{O ���8���L�����@�dR�����w���G��ʁ�j6�j�OXq�ͦ/ˎ\��Q�L��޳���md����NN���lo�#a�E� �td*�{SPv�wF}B�/a�kD{`"i4Z��,�k	�Y-�-e�x�ðC��1l˽m�w�H�gm�ƕ����Dz3��#f�(���wg{�$��=��[r���\�J�-��;��v:I�詮"�;i����p�$���X�3��L����i�d7~���<�a��eL�܍����Ǆ�����.n?!m�kJ���8՗ܭI�Ѝ=��1�Ŵw׾h�a��x�����
tB�^S��Yw��K���_ۼ���G4D9���60V����R� ��N�!<�w�QN��mZ��\�A� ��h
�!ߣz�?�8�>+>�����˸ڋ���Ϫ_i����Î3o�g#6~g)!xCR����Z i���404z憑o\T L�j��#.eH���D�.���Qt9|&j����2@=r���n�k��
<��5f<=�0��,�F��H��os�D��2<|�,EN5���M�^MI��I{Ї�?�Z�8��YG��=���y��k�Q"�z�q��E%C���.����M�le(�T�O��p�?9����D�u����;%Z4�2��'[(��v�K�)orW�h��B�q�br|�~8���G�;�v�0uS85�s;p̼�]����s�6??Q-Y��3֝%�t5���;�4;��yzY�d 3�eG�XZE�	�9���ck�(�U)���5.ᅮ��$�m�8���u�}�Z�\�d>��v�o�]����\H��~E4?z��+U�:�)Hn�� @c��1��z:�=���X�͔�:�V��e�����d��Zno ��g��5���'���7:��o�1��L�����Gv���-�o�Ζ���>>ǃ�ƱN�C�m�q���I���єHo6�w�.�9lش�Mrل["E����-Tͪ0t�o+�t�o�Φ� �\����L���6&&o��u2�0�=1eZJ=��~�M�DGdM��'�����%5l���շ��O3Dd&�z(�b�Z��MG�W���I��	Q���K�HV���S5����6�q֫y��y{C���J|�6M���>*�\mI��)5�bd�A&jA#r�iĨOD^���u�S#8�}����;I�A!���:�̼3i�@��G3�t9�0[�M�,������z�h���i���c(���F54~i9֙�Ǻ�8aԀ�ʁ�P�0:)U;�9�=]�9����9�8.O�M8���RU�W�Q�s}k*�
0�����N��p?��$1��H[����ug���Q֚�� �Mn��F��#*D�o�����*��4&��l��bs������U�n����[권"EA#
����V�Էw\��������N��}�9��ƍxL����}j2+��9!Ɋʹ��E�Ut:k�'�S���,�`��=�pL�^�UF.T���ͼ�ٌ��,��!���񻹿��/�����O�m��x"��^��@1>�{4I���U.��0Z�b�(,��s������V��Z��I�����i�۠��+���2l����aO� �,�%�2��%�g�w�*Ŏ@r����A�t�Ӣv�H�_p����;�G�c/���������wn������������I'GƳZzSH}_p���J���zXx�������1bZL躯+ZJ[<�sQ��M�����2�6`�<9�m/;
L��d�&�={`'�A�0	�Hc�;v/�ʋ�L=ڬ�\���'�:$�j�HY�.�H��H0%�2:�H�4�Wޏ!��$����W�HpA2?Uu��J�c�����Iŉ7�ӹ�^�[�)3[��5)�6!�Y�Bٖu��(��e���@�o�����a�	ᬵ�<�o�sB��'���<G�a��m�v͑#i��'�}�A���,��A�c�͛_G:�h����[؁ b�B���͢�sH�����f�;Tȳ��N쁽V��	��X��5:�j�����O!8�(9TX�w,F@�<x���{��N���/�9�{օ�'e��y�=�L1A���YwG{B�vE*M.}��悑i#J�m������p���X����5�(����+(DyԢV]��͆	�����X����(
��������K$My��)d/v��Ь���� �6�1��^k�5���0�U�d/���D!0���E]���6[m��I� \x�Y��~v���įg*C�Wg�WN÷�����8y�X���w��32�&�7��q�)\��0$����<����MVw����z�]r�(��]��B�NT߼V�G}�A7�L�Y� �3	�
�ǃ�T���������3�K4�F�ַ(��7#��:���	>O�C�'�r�Yh���0I����H�0z5
��D�>�i�M��*#��񳝳���J���/{r��cZ�W\��P�K���LYy��MI�.p�r3�-���\p�b�U65��3�|eA��*��&��/�h:M��u���@�����W,@=e��O���.�(�ɑ:�u�ϙ��"\4��%��~n�U����2��b'hW|�洃d,lg*��E�Ě�ǯ)x�V{"��3d�!ȳ!����7��%��H�ѧp%`��Cx�ɿ:j��G�w5�J{0fw��ޕ��x�����%�a��sQ  j������x��B��NZ&�.�/���kE񰰈�N�a6����G5�>��D���1$��u�
f2�±������_o
Y��*���z1��Qr���cA8Ptߴ��h����W2?������#�7Au&�����?�&�I�$��v��s�q�M�u�aZ�{c�j��B�y�X�$wQ�n��9���a�<0�f������ x�/���)�|��+�{K8��غ�v�%���"r��,����(G�R��I��:��:��ی��g|�r��͋�j��6Y�~#U(�?���[��ܒD�z�_�}��@W��2!�fz��G�\�;��\c���cr�e�r�q;��k�ط)���O����0���@m2U�ai�ix�h��^Z����͞f^��\S��w'�iqɮC��TF�a��j��'�%����`�yT#t{X�:&������W6y>&�p�5�Cy�5��u�Sy0��G�S��^��jU#g|�oE�_�ysp�f�wE��{pĉ�C!�Z��<��b��M�g����l9�{�%Pۧ~�N��dT����doH8��.���q~�G��t޸Ɍ��
��,�4b�tۓPH3X>i�&���������E���WU���J��(/�Pn���c�홮( o�-k+��y�Y�܆������Ȼc�Y�X�_���_��21|�����ȳ'"T�v�0Y9��6_rz���2E����M���%�N|��*��hv�2�x������u���N]mV��Sf1z�6a,N���l��z�e �U��1/V������'��� ����W{ŧ<{Ҋ����`I�6h�C�L�>�*\���U�QJǸM�u�[�4�ؑ�!7�p�B��h���Z�ι�p �}	o\i�:�r��;?��J7��
YWZ�r�xyS���?��Dsga��p3�a�lo��ՙ��p�13�m7�DA���V�û�W�$�ܸ��w�O-CH�K#�<��e��П>"�%�G�b�^G�f%�'�9x�͚����n(3�c4:��B��s�p��3�Շ�ifQբ;�UNy��?�X���c� �/
���[g�����J3�Xc`�,ȸ�͊w3�0�W3��AP8�g2���v���J�lc����G"�j���K����˪w����|��
��Gv��`�>jrhI���N��?Y*B�r5o�4>��:Z�Wu쎦K ���
�i:�� $WbU�'f"������5�����=��"�\��v�ƵCȑ��Cъ�H|�a��\���i: 3��`ۃ\��x�p4ٴn�%��`��S��r�D�a��р���u�֕�ִ�\�����A�5B����cv;��r��|E� x�U�x�2��: ֭�ȊP�{=L�hW]5��S���	��a}B�RR]��u��?xwV�R���q�F]� 
�D�م-�E��.<x��]�F+�gZ��kp�و�75�H)�\�u�Dd4I񬺋,���\�y�R+��u�����.�F��ҳw��]�{1� ��n+фh�p
�q^����,�t�ǌKd��*�yڿmhJ5�X���O��G�h&�C�nE7P~���O��u�_��	
��T����1��zSK�6�r2'X��ߐL�к0�T#Dܿ�u�F]8�0�?�|���y�f�"pW�D�^�(��S����==��d��!�����6t;�1pl#7���7���.�[��N���c/U��^��_m<�!��Q2�U�2岻��������� �-ݡʉ�V�Lx(�_x[S�} 9�	X��l�D\П�!��i�>V�`�Y�!������܇}F+4���DT�{�������f�zC�S�@r(��ʔ��[�H|-��2�Ȗ��ءud��_�ʣ��h�{�6c&��R��D<�(c�*/�P^�};�ݡDy(�Ĥ�����<JGVM6��%%�LSn	�շ�HC��C�!��ń:RC���+��C"Hޥ�QX	���YD=��jZ���?4M����P[�9d�Fv�)��n�K��+lDhy��W=LQ����@���Fa���)ڦ���T�ꃣ������>��ϭ%��Qdf�۾R�
v%:y08 t�S�ז���p�o��F��@�m�t�hhH#�R��y�-ԧ0\��l��\��稅N��m��3M)�����h��Q�p�a1�=�o��^ڎx"���e4��Vؚ�g3���7X-Ys�������-��A��[h����B�x�,Z�尿�&N�