XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���;�	7�}n&6/?���؉�.>����$v$l���!;����(���{mU��T��&?(ޏlWga���\��g��1�d|��R���s� ��Y���TPa�g���֡U�(��rg�t�-@o*��"f9#��߽+���9p���m���Z�/�*X��v(�3ei˹O+��/��U~�ߢka0U�A�ȁ�m0;���>1���;D�L؃�!�b�)�8��~�iB�Kx[�;2����͕K%�|q��_�Be���!�+�Ay��5��z��	�5̅벯_1��f�)�ĚpH�dN9RdV���[vI�����$�?1�x���m�ǇI�?b��v��c4z�X3��{�sG�t��6� +����cѼ���),�C�X>���V����%��-Ȅ�H;�n�b��#��9��if��%4{Ĭ��۴�?d��j璀�(�$l�)A��@� A~�{im-F��'����3sƔ�K���/N�^.E,X���m����ي���0!�_R��;6TAl�&'F9?�~�C��B2agA 9F)��'K.#9J�l���,M��p�k�s�T��c���}&���g��g����\��
�࣊�Ĕ�1��ϴ7+$^�XK��ȎFY�S����ٔ�E���"���P��n�,7sE���V�\ֱPÖU���9��ʵ�\Bq�������,*���@�&B�:#��Z��:��庻�?�ba�	�LL��2Y��FbUۓ���\fBXlxVHYEB    c763    2600�Ѻ�md����V1�CJ4z���3�" �P�Έ�~��o����#ʼVu|O�� t�"Ʀ��5���\K�uI�N�m�S�\z��ߔE(�cB�2�W<0!c�N��n9�&l�;��A����e J�o��+��i�C,	�[��E�>z��t9��O"v�G���e��i�����]����g5���T-�A����^��'�p~�Vt�ȯ�| gí왯�9�F��&ntdSN(���F�%�A@!���.���(�J9{�U�I�c��lK�ڌ*��M�����3�O=�C[�;�W���jbJ�λ��<�\�FNЦ���WUL�ݲ|�a�j%�z�3���u��6U�#���|>��`�ƀ����u�_+����Đ�4��kV{4!�izMu��o{��@s�d�7���>q�<@�%ʩ��wT�Š�dؗ���Ͷ�|��ހd�7��b�xY$�s>��W`�D����oD����y+��m;���8ق��RM2�N�����V�������A�J�B�:�S0�~U�x�E ���T�?�;�l���ŋ�2�&&RX
��MR�o�x2Y2��y�T�3fA7:b���7[i��/f���e�#�����t��|7�xi@�
�H� �lם�H�kc�/�?�̓:���EqDj�+�zõ��<��ն�^7f;l�
7:@[�=e�IE �?�TWN���|�r�j�w4�.�!��l����v�����.T����I�7Y�pћ B��)���
�BB#�?��Ax��7�mƽ���hh��ߥ�{���a5[
\Lܑ�K��ɄYŋ��N�3�� ��1��e���Z��*{����S`�b׏�o}Rl���4���� ,���[��~6��E�,�ݎ�a�ڱT��H���K�z�}����P�3ܦ&4y5�7>L$��������/k�q��oa-L�zs�M���ҷ��m��֍��e1�2���F���L���c�M���`Z�O�lX���q*>Ã���U�"ï�Ŝp��H& � �[0�iYY�h۟�&�H�~ޮDK��'���@F<�U�u�A�'ޔy�m�i A�������Q��-����&���	�{/؃�㸊�8(3�il���K�W�(���=��,v��Gv�Mz�+�H��	6���-���`Zk���Cs��w�M�b�\Yt��-�|�y�,r�	,EGsϹ�5��
��?Q��!�21�z'��)M��h͢H����	C�fr"ş����_�W��(���Q�Xɧ�[,& � �׺��u�Q�\C��1Ip@�.=��d"�B�W���^'��t�>Y����/���ԩ~�[1k,L������#�S�:T�K|[��P/��pN��#1tȫ�4�3Q�����M:�g�Vy������Uf�UVfF,O�F��������;/*��rW�qz��c\�����k\�n�O#��v.!�/�q5���筚�o
�Z�g]Ψ g�e��Kb��>4��>.�n:+�%��7��-�3�e4��m���X ���gd�m[\��������Iu�h���qKɒ��O3�k3��<D�j	�Ra�F�Ϳ��L~���X��3 �hL93{(�S&; �l����mҔ��eݨ�W��)�>�$��I,�|s��=�C+���&�#��k�-tZ�Ā��;l�F��V���Bæ`��Zi-ש���Yp4Ǹh��\��HƆ��w�7��Dܸͦr)%��3Am)Ts_��x\��fq���.����dn��Ѵ�
HQԚ��.����N���ϋ$j�p��a��]zWݻ���gdP�΃��7gc	��e
�	Rw�w(�U+»�dhh��Q��d؛94d����%jȌ�֦?۬����`B
�����4�?�p	z��#�?y�`�"lQ{dH�$�9"~?f�~�gT�E��~X�z�2+����z��W���L�����1�q䥹�`h���`�2uSǑ���U�q�t�+ߐ�Y���q�2	g20l��Q�9�ηj�UdK�5턹אz~]�<Z;Zbf�[�B��	Ƀ���덪�cc�ŉIBǧ�Kl��O�ʾ�v��X���;�}�"*A��$�$y$��J_5��.��|�IwQnԘd���՞�g������)
�QQ6U��:A��	��O��b��]	 3$J�ե-WUX�1�����m��4�~[��jӫ���d��k⸬���V��S�X�ţ�y�h7�?M���y`J���H`ǜt��{�'=�#�2���9�3�mh~َ1�ܛp!�hb����5��&�i��VH��i5��]t��r���-��p��ډL�BtQ �z��rÄ~>�S~6��p�6�КlX�^sO������[^�v���=��q�px��j��_�[u�q�|.�r5H,��`�R/��=yʑp�s��,���Vղtͨ )2�u��]Y1��}�=�-/��^�sY$�l��q	h��lӓ-�����s��$/ԍ.���ܟ�Ns�U����MִЎl/HY\Z�Y1y���R?N�J����C}%�B�~:#X��P:f�MD��oS tE�F-YŌ˸��ls`��j������0쥐�L3��F�ʂf@xϞ��람�x(]fc0���	Z4��ԇ
ӆ��n�P�q�j��f�e�\\MI��G��n��ǎ�?t��2�����I����2��`|����2["��25�a�"'�}�k��@K�y�vcV���{#�V�Meyd�_���-N:ѷ�-]3o`ۃPd�`���`��(;.kstP����s4g�{�6Ӹl`%m�s���ý;������=���r�;	�s&|sP����ݔ]dQ'@��嗔`��H���n�x�WK���x��Y�pk�X�*=�Zi�FiW�T��Z��ok�+v��T�y9'rK��׹��g����ʏ����rT"H��� U!����3���S�Vv�Sպs�1��Ga�}Bu9!<���}3���m]ʄy��D�a���Ò�߀���BA˺Fa�D�V�x��k���� h�Q��y<й���������9zo���p�|qڿ��k���ߜ'������=�¶j�}j���������5);q�~@�|uOPv�hF&�t�Xǜϑ0��+�)*,��&`�s6�2�#�3�t�=S�5K �2+�Ņ��W�^��Qn��df�"�o���ףz��%3��9�bKW�Aՠ�B�>���]0bF)rRY�d��AU�X��He_7�1|�w-D��19Ap��h����a��9 �o;]i���goB��.^i�Z<2+ԏ�������?Z�
W�-�k{�#�9fk@:6J�
:��֎�k;�.�Ha{+���2ZoO�U��/D�w��w9�Qp�I�BL���ʗ���5���e��O�'��+�xޫ=ڄr��/r�;1v�2��8��h5KH2�e�A�o�e�*<�v�w� <�q-��j�=y庢�&[����X���H���"Ax�?��i��0�;�����[�C�M��keZ�P���n�z�TΌ�R�v�Vb�R$=���H2�9�/��]��*Ѵ�b�2S�<90k4�]�07����x��0�<���̟hXR�Bdt�|��N����Y#	
��E�Oճ������z�V�n�U"��&��\J�ؠ������C��HT��RL�Qm��B.��3
V�����}��fV���=��
^HKzX���2���=��t�u���,��)��6��N.*5��I:rCB�+��67�东��S�
=����xO0?�^�=j���LfC���=n�4��:��hG��gpWM!���M=�ԼC�#� �m2���9S��t��*�������HN.9V�ʘӕ��o����l�l��%����0�[ݽg3K�ܪ�Z<Ca�~��,������z�Bu�q(��qC�����'����/ِ����ѣ�%�z����oB�ϰ���X*�6��H*���ߙ~4���ZZ�x�gS�ǌl� ���&�@�d�2�*�Įzg��[yedLQ*nK$8�J"^�6m(���t=�5v*"�nV� �piQ�-�c�-a�8��,��iF����aգ�qs͙������bm�R�[0�l����:D�XhHn�uS����W`��b_߇R�M9yޘ�_��N�"Yq�b'��p�Ɨ��k��{լ�l-�/�]D+�6/\���U��6d�@�h~�b��LD�K8�hc��ś2�mX|B�{i���[B036���z�[��i��3Gт���F������-��Z#�0��k~�~O���'J�T'�P��bt;5�"8��cΓ�!oc.'�	������I�P�����]t�������lN<�=<�j��xMM�?�;	q�����붥����QR�x����Q�jE���ۛ�'���X���Z�ոU�(�bk��. W�|A-��g��J:�8��w3):��7�-�9R��Jd�,���ۻ=R�	���{�$�ɜ�gBs�[65ZS�M]G�壁͟������1}�R�	cq��ެ��O�����w���\ѳ�u�_[�_~bU
��4=6� ����������Ӧ\Vۃ���
��V��<~�s��ʾ{	��_���m}IhYò{키�������2?OU~V�1���;>�=�X!|Y"]?���4�W�����/(�ɭ}@ap��	�[̫ø�� �����/�-_���HβNv]J���~�2M���ބ��+7Gx�0�q�g��n�]�:SN�>�F���h|d+v�O��{��=.A+*��������c@�]�vL
u�(J6#w���������ҝ�[O��A��`F�	�����09r����B��XI�2�����7�Q�����zpvv�ug��E"��Ĭy�q���k�lHzzZ}���M5cM�o��L\�,���L$���2 }^@:�s�%�h];z|QS'�@9��\}u*����(�~�!��F���)����ygz�|�$3�[��е�r{�ٯ���`4�9O��s�������߿0-(ۃ
.�� ��"ם�*�:�Y�y֛�p��sRbG�-�wY[ �����,pw��0VF��lL�`�����r�A�T���L�7xs�O����C���@���;8U�<N ���K����~R��2hXk��n����+Dk�	Z��]Wʹ@�En�;d<�c�|h �&�ݶ"��pk�[�4-�a弉��z���{sj�J�f%���(qb�%�#�?��
@8��!r<�� �#'҂&�u1Rj����k�-�2��}}���r�N��(1mM�f,�j\�gV6r����7f~&ǌ��������	}Ja�����?�p�~�ޫe*��`��&Ed߬��Bء�g;�D����ר���v*k��,��Fj��.ؔ�r([�tPA���{>��"9b�����:4��䞬�+�Ky���/�.o0��-
'���d� B�և'\��C+{�����"����x��*�@u\�+7�^&����vzR��t[��MAnm���ˈ���+�����ˣ���;л���f�X��q��<}2��� ��g�T�K�
�gb^L�����/zO�S�tn'U��	
9/��:�h�O[�b�H,��mB�>|���B�L�O��2�O(P��)T�?�{����������z��`�e%�ʸ�JS]㧂H���~�G�w�k��ZZFl�\k��
��=���]L�;��]@H迡=&���o������(�;̆��b2u�>z�X��og��w�����2�����~Y}���6�UY�N^F*��N-W2�U��U�-��.�	���X:�Zz"���H��M�ҕ�
�׉K����{����\Eh��`i-jiBg�5%֝���W�x(�R���	HD�;'V%S��d*5�ҷA���LZ5hӞG�mt&;<�^�S�F$���g�*�I�#'��5n����c~��&�84j����K4��tmly�ӟ@�ǥ��!����3��;+�- 0P՚ϡV�m��໖J�� �c���C� �k��#��*�z)���)��2ňhFBK1��0W�?���z,�5�پ�� 2p�S�.��kE��y��5�'�g�j�����dE*���kl��߾�	fZ�	�L*.s0`��t���sp��W���z�7�[�m2�^fr�Mʻ�$ u\T�E!<���J�����2A��m�^��N�b�ʙ����k��o|��<Aa�|G�m�׫��p�)R�ֱ���
���~��d1�����z[)ekr!?����7G�g�S���u R}����{G�������j{�o�t�!�#w��p{-x�xㇰ���d�X�Ůe���D"��I�� �)Eh�q/$�oc�X_����Ċ9T]~(0]"i=��K�SV��v�e��բg��E��d𾏾����QZ��PI]5�l\��y�p�u����9�hڣ��2��F�bm���C�ܥL��8gg"����!к�`K4
-���H=F~a�,F�r�ߏXZf�pAϑ��[`l�|��	�)y���uE)z$���L�8Y1{|��^��䱘�ܒP���q�9dT|�0ϟё���o��ƕ��
6ʳ��D.��O�7���4�ߋ���;�~���Q޷l>Mk�=���soV��CJ�K�	:ԁ9�`7T�x4ađ�%SP5�T�|)�R��L���ޥB����m����G�2]Y��8��x�fEY86E���l<�T��c�쏔�T>�m�
�T�M���J����x7�!*c9��%�!e,���:�|��\�v�����H��P?����l��8��"oFǱ�D6���Nt������#~ؿv�<0��~���jk�������9Qځ���jԒ�v�o����;��@�nz��v���}%M���X@�ahK��[�����
����9���	g���W��$mT8� '�A|���rd#}ݾ�� ����8�q$�l��O�â�	��U�T�P6KC
|���š|�hgl��6�y�j�����.�2c��h�;�#ě�5�f"� �g�g{� ׉�
NGH�����2�Ŗ<������&���7�FʑkX�&���_y��SLxEչ_�����Ͷ��!�:T4�Z�R�!9: 1&��;���m��+͚H�]!�@��&-��s8�&�m�����^�?��T�݇���������p��������*�Z�98����G���?!Cv�ccaQ�O_��~Y7�ռ���Ch�h#nh�T[�����{���L�v}-и�G�\��������l�c�N/�8%�CJێ��l�@���Mn!.&�=�
���O&Y�m}�d�Z���0�C5�y-fF�\��JZ��]*�F���{�ى���?�*b�F|a���%8eszn�z����wg ������n�pQ�N���:'�w
��y^��N���r#�eY�i������ﶎ�y/l���:����P��:N�j. ����B��;Zҩ�a#fB"�T~n�AEe�H��+���y3��%��a<(i�k7�ST���
��c�m{�����8�����fj9W�a�\I�V���,�T-����Q�1�ɢ+ֹ E߼�L���v�"%A��H��&6H��F��,�_~T��i�L���w��#Z�A�F����y�U�y]���h��x?h)F�����ӧќVLٸ&!EUnb�98������	� �y�#^�Aϖ�����^�iK�%�V����m����t���:2�no�:�V�k��%d�sy�N���N���0��	v�Ս)����d0r6a�F=I�sf��l��x�k��V�{� �ݶ�u1�	ՠ��H�1�:�*���u.G�#�O�d��� {Αr�	���K�Q7Mz�(����?}�����[���>d�jc=x���q���Z7v���yԝ�+�i�ˮ�򲻿���v}w񏟨��\\�ش�^�@$?��vޣ[��"%^cSPD� ��KyK��?f|�TW�V�r/�LN��.N�]@B�}��񈖋�W�Ld��y�\�#:�g��]��h�l�Z�
��I�:����8uc9��q�f,�6�Ƒ�b�f�g���]|0)i�`gB>�+@�,�%N�@ z =���mys"�*g8�g���vY*�,��5v�����a��G^_Qi�<C�4�^�=)(JO�ʢG�����D�����!GY�4Ӕ}8��	rK��a)�f�b�U�qo_�����a��8*�u41���WZ�J�2��}�Ly��YIC�E��,��'�.=�U��m�h���e�
�2j8%�s��Ue�����0z�r����1�&t�<��cd�h�+
+���aHI5f2e��~�i��cd���=#I����Pg���q6�p��D�,�J�_Ex�Z9�J"���^~��/˭�p���������?.M�M�S��[�%��*-��G�b@�� �R
b\���9��R��������BM�,���pށ�|����d,��c'���-�GXJO���9���͇aFMS'�!,��Yz����p��<A���51o ��6�����b��K���|��I�����E���"����cnR;D=9U5l^�CUTr�pN���g���O��˅�5��8��%����j��	���Κ�K�)I�t��R���4�-�N���t9����m^ �Ŝ�����ύ|3����\T}��`g�K��;l:�Ҿ���:"�����I�j}9+�Ϭ��^&�+W`LkR�c�}�+�� F���_?���=�3�,�n�(�(h��[��0���@,*\0Aŉ��]�v����n�^%����$�z�kW�ҧ�gN�VH2�5�y?���S�5�"&�s0�N�H��9c�����]? 5�Bͱ	G��l�l����ϊX^�L ���������� G�g���o���;�Hq�&���A�Ϥ��!�n��_�BO���s�+�F����fʗ�ͼ�P��Fᘗ(S��f7bK�^IfsS@;�D�Sk4\>o(��?��g$W�0� �i�R�0�Z�Ls�xQ����s�$����B��|pg��u��D��������v�����1B�vIfq�mn[��
+h�ȩ�Nr��˫Z����ec�� �(4p)��Rc��Og����r��f��CCYn�����+��_n�``�~��8|	�9�G@���V��lg��h�{3!���}֊Hȹ>�\�5�R&W�h ���*�[x}�hӶ��r���@��{�YK�
:�C�4�Ӛ�3���3�S���_$v@�J�c��_��G��c!���$�2�����M��D��{(����z��q�!��|�%j���H,s��@��Qˎ(`Y�@�ׅ�D�^D1���0����`��w��5���QSM�E�s$�z��s�zл�%+��յ�]t�ڦA���eN�p