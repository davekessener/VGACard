XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8ZT,f}�1���m�c�6/�](�TS�,ԅ��,���S0��`Ģ�o��j&ڹ��;X=�?�*&]��%��e��Tr��Bv~�|U����-����bw^����g��+��ב+���'�ߣ�P?�v��LJU����o�zFA*:s��㧠�<^������iD/���w�H�~ ����!�T`o/O�!���[�;���5F���P�>�bv��.�o��xR�W����p82�o���-��`SQ8n�o:�F�d�`W�c��(`j�i�ף�);x����f��O,��㥭�'Zu� (Sm�L��B���d����j�)Z��:g�_g��~S#��5%��L�tp�2(���Tg����b>�~�ķ(����Bq����*C��||�J?�%��9��F%�H�ȡ���4����!�)c��E������v�h�������9źǱ�~*��!,yu����P���7�.�M��z^S�?�<�!s�=�����-�n���Bt���O�Sv`�3�VW�}y���W�)م_)�Ճ�U\�\��M�<ˉh{�� t�(��@�7�q��C[�k�Gtٙb6'�|�j��(k�r�~TJ��*�(��k�-a+�������Q��m�����+��n5X�ȶ���O����yJ�(3�M\$��O��]�B�= .K��*��O��UG}�S�-��Y+��k'�ˮU��6 %�T��~�����1��<�H�!�#����3���4s�T�]������o���njPn�?XlxVHYEB    1427     840�x�+�#)�&�▿�A��j!t��?h�U<D���k�` ��3��P`�pcJI���s���� ��_�r�.��5��,쒜j��c���G�rY�A��O"aW�S�(�!��`lC�4n�X�ǍC�)"C�5<N8+�]�;i\岦������'����2���?��D������d3�%D�� �1<�/Q�*q�*1�&b�e���8,���ἳO��6]e���F�����A?�w���/N�W+�؅����~��X�AQO"1�L��$�Q��n���I
��v_�4%d���,
�.��^D%�1�������^1Uf:(5}v���[�'��\ ����^�}h��϶�`��Z��'uz3�~�ؗ@�l'aPk��`��J\b�w��J�1��<Ě ��ZoJy�h?�y�4�n�A�<-� D�?=�v	�o�[�YT�GA�S��n�r�@c�h�%d���,9������ca�����8Y�s� �kRch��4�ќ��t��W��ȳv;@z0E
)����:���>ވ�7�
7+�ek	�KeZ�W�X��z�_k��M��+�M�����6?,��M^��I�����d�!�YO���5h�<6��?P
g��Q��*�h'�6uݏ	9�V��OF�a��!&���c�l���ͷ<��1�}+(Jj��r���~^�"��{u���ݸ��&Hۭ�wL�&Q�VT�,�a�Kz��E_������Ct�d⨄C%�0y�� I�^���A�R:ɪS�-\���w�B��R���°~;{{�D�Dw�Z����7�ˮ��U��b�v�7����#7��e�X���m@�ޫ��ں������
}	�Q���d%�|�����cmB���@L�l�'��L����f�Q�������ɕ�{iw�K�Pb)�d���]���ف�-�%��E ��>(�h��o�t�>}~r���Ն��t/�n���x�}Y���R�@�`X�K�����{��iu���+4������q�;t^@r^��E�]j΍��f.<�A��>J	ɍ5�T�^�Iٔ �l̀%R<9n�Z�^������8IA���{����Q{�ɕ�&1[��3*��S[��$�\�L�@�ia��}��"�*����(��A�+��|���n�5�ZL��M�%ʲ
4���|�(xV�uIM�on����R"=�H.���]D2��~�1f����p]	����S��0Z�e,�6(/	k�v�(���cx��.N(y�9km��Ph"\��4v�! ����}b�LR� ϸ�k�l���ѡ�H���Ŀ�Ϧ���V̓3:G��Ȃ���@p0�!uA�!Ñ{��Ve���&�~P~�:�c��}�R�N��-h|"�{Cu��J������#�����:E:4O` �)�8�Gᾋ�����N~�S���M��g�~9T�5�&Y^��4�((#��׻1�]�]�w�JI�2\��<P���#�V�3�V�Rt�E)!��J�ַ��:.�ѿ�u�"0Bp`�+0(�t��|�գ�=EYA�&74R��]��GbO��6m��7�|��d^������#���o�)�S��-f�W:���Y�X�q�1=�!M\�h3�˳g�ߊ��'3�̡O�����\�����U��G��_�v��|^�̸d�2�?��8Z��8b�CO�¨3~6��x��d��|	��}b݁�"�6,�G{��p���TLf�!�KvXm��v�*.^��ם�0<-��]���$��_2��9���������"B*SkI�^�8uŰ:�Y=��X���4<��G �V��-��s��d�Z~h�Þ�e h	j���蘎.�v���u�v��}*����߮#H�a�K�̤jaO̙��`g��fy_���~F}_�a�b������sbStxN�p_+���?��]�ծ9�6��G;�4��l�o�H��vJ==K�R�6n�g=�������UꝹ �gʳ�T	�V	��b(�J^���}Y��>1�8F�Omz�F��^�lDU��U�b�=����� V'윫T]b�6C��������