XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ce/(��uI�&��[<,�����_��$Wr*�U-��W�+����E�[�D&���I��.ˤ�f��b/
��&��9���@ٽ$�S"^�a� nߵ:D#/���rQ�/�jv�84�J���	��M����p=(���!�w���B���"������U��uO��K��D�����G��W�9iUe]j�BX3;�A낖 ��`	;��6��V�z>x�رZ$���M�L���A�4	�讧|��c)���-���P��lA>h�0�9�R{?/�I�)t����cل�j�S�����x`O ��$�Xt+�lt�F�[�
�^J���N".Lw��-q.l<�X�?�ﺜq؁�=l!�X<-4v�u"�/�r��yie>xh-������p�W�[m�EQh���:��\>���{��%}D;8X��Ah�w������"�
�`� �Vq4�~�%��@�|�w�T�IR�r ����"�+��N1cf�U����7� ��J־�4���L��0�5
%�*��P�0�W���Hbլ�J,-��fe���2L��UZ�� �\�Q]�D���3?�VL�O�h��r�$-���þ��,�{���zӗ&�e]�k�B1���r�b�?��vz�nXEr~�ȳ��(-�?Pd����C�������q���ů�R0�ƄXie��pCK�+ߊ;@	��i`�����<�צ����!���m�G῟�q���7�j�85���b��m�;.� V�~XlxVHYEB    56d2    12a0���u��3w��,J���K2Ji���v��SN�r�U�w�����= n�S�:m��<E}�����Ta�1���A�Y�kA����7U�.�Ϧ۲t -��Q9�3����������� I����P��b�b;������v�*2Nr O2�/n$gIR��c�	g4���VL�W7n�P�ܲN� �L)US��̇��`=���^�%g�1���3k�/��σ���Y����n��ׄ� �ټ��PFwr�;�JMk��کչ�L�}Ũǟ��Q-fb-���,$V��X|�n������3��M��_�(1�=�+�V�)��^b��w�x�u�p���T��"�ބ�ȖI�Z���c�����Ț�!��a(ȓ���)G'����aʠ�תO�3)�,]舎�n:�}uSa����D�!�o��`q@0�Mf)�E�n�h�[��/y��;���\��S����ϳ4*��#�V����&G�z��fJ������.}�h��J�M|	��j����e'�H�5������o�D��/5>X3��gK��U,H��ݛsH>z_>U���h:	����8�=C�'�RʁȻ�H5/��$�X��5���a������ȑ���n��=�������b��K31����2�7o4�W5KFfyTp�Q-����%K6i��tU��nJgAR���U=B�hz�a"'e�U�:����9c]` E$@�����l@��1ӭ2�ͭ!Ɍ�AeS_��RqeE�0�P�NK"�މ��|B�u&19v ׂĉ�'Y;d�NY���C'�D�P��Kzh,��\�<�Z���BM3e��b
�C��s�P|	�ȺE.͊Mk��	����vł�#+�U4�8*F��0�+m�i���<�_{a�)g�ι�����]�w7�J�bx'�l���E���J��#�m�m7"2ơ)V/Ý���<�>JaďhG��a.�#���}^#@�Uv�R�5'֞� �D&O��'@L�!]؁�T7f�䐭c��)�[�,�
Y2�(�z���6߷t\��S�2��B&�Vb'���w���+��KzX�_�\��i����g1�i膂��ި��>�N�{�Z��d21ה��_>��޲���p���C8�]h��[]��8�� ���1�i1��\@Q��0ǐ/��ܧ�o"A�5b�Q�0ɏH>�hYY�窀Sy{��	vL����ι�w?��j�A)���BRmK��_Y�9�w�)���l�����@#�����q1>4s�(���13C� �ף�QA�j;z����NNj�J�n��A�l]/8f�L0�l��c��<gjd��Ŏ����sF��
�T#�#����^ym�ZDj�����6[눞�q�Z�-���H�Z�$���}�_p�$����I4��Kn��Nۑ�J�-�vgr��,;��:֕��ƫ���By�yh�`����f�GQp=�Rn���$D�2�Ţq�o��1FD��l3}�Ȃ�p�$��+~S@H�	�.!�2'��سpq4�*��Ƀ�=��GY�������/�l�FG�� ��o^�:�!qwk�P_���b>2��.��<o$��:�f�ψ} �I.q}��ʣ!���`O��q�F�!z�f=�Q��AR�/�w)d�pw�r'c�"�G"�X�@���~�`�)+�c֧��hM�ך��-�@bZc�wr�7��z01�/�ȹ%��&F_}i.��E+�(�j)�l��R#�(�����M+0�k�'ۦ���t�3H��X\��ԩo�)�ײ⨏荖����c�D�yn��:��s^|�V�#�L�hFR>����꾄�긻��h4�:���`���Խ��t��Jrr,
�?Hy<���f�M�I���2��&�=m�9��2a����FH#�
�d]x�\^r�H��\��2Ѐu��cc7Tm�	����>��ʁk'�?�"�,ک�g��&�wOCx� ���������D�"F�yd��5�x��.���pS�RS^��n��J���Y�R���7[�u 멚��v��H ��"݈=Mz�7�wS���b��T�i@^2$��
�Ք�������&vkw���S�+�B�C�F#=�(�v��G�g�·b��� �0:��Zp�r�@��h8OU�( �ΓG�k�� [����co�4U�9F�o)cn�F|��O��:"�V��	�7�y�/F�깨�g��>�z48�㦐��5�9˕+#Wٌ�������9�d� ��:����1�h�&oS�,���ȁ�!�����ᘗ� Ά�ɿdz*^N`S��"E/A��DrIGZ���Q̶��'[�~_�Y�W��U���!�����Һ��
�'Q���Φ��e�1��z�m����m���:���g��Q��9H+���`!����iT�sx<!Tʮ;
4Rtݫ�	��D�ә/�ak�?Q�J/T!qz~o�ku�[%U��)5�3�)�RNn,#V�}wm<��J�B��w8C��-�9�f�U2Uv�r'���s�|��*}9��	��ZPϿ��3@�qE����X���z����n�Y�´z�[&��>(y�2�=�����A%��UB�E�i��y�7A[��p���@�n�V��n!=(=��]1RS�z�9���e�����K?۞G2B���_痤����o�~��/SS�1<�K�o�h�2U;���y��6U-8L�w�fZ_>x<4TO镐�OPKJ�.1�(#���f�m+��aUI3�mW�	:��Ԍ�����O��o�D��n�����"t �*!���%g�~�v�4i_͖0���i�4R��#}K#���!	y�*X2��Q5ԭW�5Y�|�Ku��M;��ª�m�k"��24�/L^T�:6��gt��UL�E�-Wt"3a8G�!7���5��􋇕���`$[����l*��r�a!+�?��'�*Q�����1~i����V�,��@�����SR�J��4�R���9�v��i���e�嶻�+5����Vs6�i�ę�d.(#��Mb��z0��w{�MT������y�Ӈ�0��ɘw�t�t��0�r&�ŧ��/C�T�w<("[�s�{񈋦��!�v��,g|�z��!~���"�b��f�^�p���!�y���ܽ��-�Q�7��,q:&FR�|F蟏w���BR/�3) -�6�N�s�]�=�GHf���w�3�A�޺�h��ur;�!CWu"	����a�&�UGȡ=�zQ֬��Z�bu��&}y�X�p7[E-�x����psʂ����-�26f_EK�u��1(������S<�fj7��&��k9��v�j#ť@��z+��䗺�FL�I�QN�ف����=U�3|&��A�\�'ԋ�H�����%��81��"�a'�'����S['��c�23ݽ�aUax:�m-M�#���~x�l��Ym�6��+��I��
_W�8 �S����S�����ӝ#%���eN�8��-�3־r�Oy�2�$h��hkwT�`�U���sG�:)��)�Vm���*oH�aݔ,�^��j����8���{K�m��]�p�Iܜ��1J!�}�0�FP�领���Ƅ"�=}ylǮ:i�&�;)���Wǝ��B`��s���l�CU�N������o��Ҁ��3�JKy��	IJ��2)m��舋��KG,�y�U���=^�v����)�X~Żd;�z�X�ɝ����0�?i����3S#�������ծ�;N�k��cwk����k���A���Ѫ'�eS���oPb�R�Z��� �4��$I���{)�q�$�ر��a�
��1�1W ��F(�X��BQ��e$�%�ҩӕ'9��K=�y��4���-9�_#���'�Qj�x���$��H}ɵ�0�H�o�w~��̵��O���^SN/$(
T��U{~��?���kOM8\�+���w��}���wh������/�0r���Z���x�#k��0���sy��cy����O�e�)���]�Nu�LY`�L5W&���p؅A����'t�6Q�f�� �|J�b2#�l���[�NRq�S�Qk�� ��C���<�4�+b�#����-0��NB|��}�h�T&���l��!+��J�\4^�s��5%����^ C���I�-	Bכ��R��9�`Ȳ
��Uph�́�%M?0^�3|�f�u:�`4%����&R]jA8�s��Z����,L#5�	�B�bO�s%-�E����UΖ��od�%����*5�cC~�e	b'�O��f��iĀ���*I3�9b���k�_��
��lFe ����^^"�;I��Td�5�����*�9�jھ��Y�.㍹�y�%��%y	D�~��R��,'.ԉ��'��ǘ�! v���.��8���^��mԴ̡�S���Kg�/T�`�m������.�U_���m�h���h�gj����Nӝ�;��2��_���^�"<����U|���{�A��9o�1u�m�I��KiA~#����7M�󕏩�]t��x�ks��ny4Ѡ3}��ۙ.� @�Uz�'?&,�v�"�����W}�j�R���&����w����H�h׭���>�!�I��hh��Mu8r�"(sݶ��>t*��C��g��S'��5b[�E����g�*p]��#s_P���&���<�`�Q�ޚ����(`�=c��4U��ϐ.y�