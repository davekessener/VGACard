XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���c�8�BS��\�)��`h3�!ȯD�r{�<V�=�m�C��2�-k�ڗ���� �~��%�z����cy?٫��N��[�b�3�L^o�|4�C�%�������c�E?o��~������q�!��e��B�g����p���TV�`����x�^��<�z��
?��\n��U6�����]vh8��8���'�t�}��<UpP��Q�I_	x?k�~`�N�2H����:��~F�F�
�q�Lkc��\><�7�4lC�����M{N�AtLM�UOʲZ{.���>0�kF����fSzOTj�e�;�뾼4����m}�~�Z!!�eF�+�|n(@I�Ȃ:Z1Z+���]�T�k�ލ�g���Vu���o�ge�������=�;�(��>�L�(yc�j�dy�9:��`[`>��'������~~��sa\D�b���40����5��lY�Y(���2�pk�	�&�_��T�6�zJ� �>�w�>��ޮ ��'M��ܻI�%-I���j���M���3핓ʹ߄3�<K]m��&��[�F-#A�.�]({���>��N���F�6h�ځ��^��Xm���{��4�/�  ʯg��!�(�+l�~v���Ϣ<���ƨw��7�hb��`U�ʸ�3��C}2;��k��cq�1�J������QI��Jv��Ο���,#�;sM���f��EА���q�W9=J�%ZԐt�r�T��*�y��mB�u���C���}r�2b.����f�~&�XlxVHYEB    ea93    1880I��T�G۹[���V����&�Si�Φe�a�"��1�X��
_IRU�R��ɹ�`x5����j�!�PE���mbP�!Nۏ_E���vR}"�1fu*����g_q6�6 ���t�~�����P !/]]5^��5D����S\��MG����%k�a�6h9&��W��>SU�x�O�:��Uf�H��!L�N?��UmG�3�pjѦ��?���M���nɎ����]d��K>90�ʎ�"�.� ���6�\j�˖<4�H����O~�	c�o��S��_W��'�1t������pju�!m7v��2�Eb��9d0c�#����s��}���O�\EΉ���v �3�-��$�fCS�5=��_F�9 #D���[P^,lu<��\����(K��2Fi�O����Oz�����C<dXanA��o�\�o���
�%=�Nn\�m^]�ٙ����Y��'��N@�20��>�	��Y?�.F����(Ql�q�ozNӫ�9�7QL
��<"\hfE�m��Wo���d]>t��dj3�*�(�e�;��"���	:�hF[7t,�nqwХ�3�k��^Z������f�^�aP�����=�A-��ө�cV����d�go��t1��;������2D��
yMSr��/���2�8Ƀ�`]��z��FA�^'ݩ�� ,��5��F��HT��U���ϗ��z��"DA>/ꐖ���8@)Ku��]��M���M�w�_s	�e>]m��w�05��_u_H�����.�?RX��O�7E�974��tf�w&�%��*��bBzj�Rz��$M��p@�:�ƓV 炚<q�@f���Klx�ͨ�y��Ƚ��jx5�``��21 ��a?���K��􃂾$�^��Pӡ=���4^=�Y���$R�Jp��vX��{��^�j/�����n��׏��׽΄M� K�(�E�]o��V�ͨ��>� 
�Zj#c�W���n���6�=�?���t�;㓒z�3s#��)���~l��݉(��G�9p��W|�F�W0�ؗ�oAw0N�dЍKq76E1�	a<�g�H^��M���솥�XTD_84���������&L��K�V5x�rƼK,��F��$d�v������~�b0���F�'Z��	��h��I�V�-eE^��D��X�o�S�|>�C��5�@�A�ޔ$u��Pz��B�S�0��ʐ���saȰ��n�V��+���,�ŇraЊW��,*��y�!{1�DW�,��G�n� �	�i	Q�J=����u/�6��=�>�\T{%��<��e��M���٢�������l)���DOv�zb_ �K'e������(������2��-(7��D���Cgor x�;����$����	����E�W��u�K�/��4u��Huc�3���Hc��8����p�98'w��*����������;��Ά�%��,o���M��0s�%��v�.�Y��5��p��6	������ϳ�������	U`>��s�<Nj%������~�����q�[(��!������h�~�<�Tɖ38:���,���Цi2s��^b���^'��2�^d�W��Qt�%�У��皉*�t�F9)h���$k��$.�]9�%�Q^O:}|3k�JN�s~.�k�C��/�����_�����s�����0������`�7c��oV=��J���3@�;yN.���~����򝚬�f��I�m�1"�� %U푋DO���=��t5.�Nu��t\K%!���"�8�����h8�b=��9\.�+��t��iB+O��x�����u����8���� X�e�P��A6p]���[�	��z�^N�*ҿ~�y4^I�0kbV�

�r���p�A��>H�sjw-KXr>n#U%���`l���o^���G�����)v1�^�7�I���B�݊[�i�q���e{[f e|� ���l�VNQ#k��z8x�QU��Dֵ�"ߺ�^�#i�&�i@��2Vdε�8��N�؎O�4���;M��}���M$�a���\`jo�v��7?�ؓ��4�K+�]6�e?�����-@��t�^V�������8P��c�H�����,ͧ�2bX����ZU�����������+����p+������������D*�� UE3��Z��S�� �0b�����N��ԓцa���
��7�Jy-�������xs|����-Ɔ+ܘ�X�S���ωWE_�օ2/P��6Kk��ο� �K*��c��G�'��-������\Z�yw^ւ'n�!�*::�Ga,��l��׋"L�|��1��Ad��V�+XWV�cN�8����Y�<T�h�2�
.�Ʌ��s�J#į�NFܙLJ����Ϗ(��g��m�(��W
��=�Hٍ�IY�����o�����XQ�C�"�@�����vq����_|��B)� eD����sE�*��79��j�H�N�z�U���|y"���%e������s�Ć����o.�W��Ė����~�=wk�I/�!/b��<����d^���<�%��'g�0+��=1���0�H��͍l��Ӆ8��cH�0���b<��Y¦�+�bZ�a3�+�ǝ����TiF�Tg�����vw�� �P	ep�f�\'2Sش��9a/�`#�l�T��<ǖ
�������(���H6��{�(!,��rK��a�s&]�K�i��n��[\�q�U��X,� ڻ�Brv�z(�Cڭڬ"��>G�\��>Z�OЩL�
�V��F� Y!T��(č�������H"$�)\�����g����n�m�w�6_m"�ݔ� �/��@��z������f�8�W�~���ĉS�f/%�KNDǿrtc��ٌ�2��t����R�T�.+����	Ɯ�@��1e��ڪ+� �e~ڙ���R���>dt4)���֟*�вD#x���6�����w9J"){U�y��(K�+p��h�ǼY�Yg�6��~�n{!W ��>8jX�{�M��+p�ZNR�?��Pr��Mk%�y6Ǵ�`�mT+�%�c��y�S�1�3�o���f���b�(�.a��3e���S7u�W��9�#/�V`���ߡ�d�1����=Ι�4CU5^��m�EнC�2�~I0����W���p/�P�_�S�(*,]>����r ��	<�iF>�;�;FR knF8%Õ������3<�Q�4��r���> ���F���(����d����xu������A&�k�l7zt�,�-����,�G$t��E'��
�Խ�}�̄��b\o�Z�QЂ�^������דU���Z��sd{��f����d/q;�
����N�]HV }s7{�c1C�=`!� *��л-ޡV��0�G����<��0��z���ƿ��!��`���)����G���C����1���O<���INt�n�@��a�e�]9�L��oGM.
�><m���lL���x��9�]t:����u�ŀd�f���ׇ��6���.������<���@R�ՠPx"W9醡A��c�ND]�8�;��ډ��ׅ���j`�L4�``�4.����Ϸ��x�+~d��
�K[�A��CM���=�OB|��{
o������8���%�֒{��I�:هF�@�����O�H��Wb��#?E	�0 GF8���C�F�@�+@� �ۢ�
��υ��
Q0��Z�CVң��Pv�Ee \XDA.�����)�wQ�%P�`�\;r\0�/ 	�
�$��u�����'ˑ�[̿U�ny?�_V*�Q#KCX�OS���"�����T��we���4���TúT��������2	?CE�����y]���vd��*�p,[��X��i�#2��P$䓆`8[lG͆>�O8��w�q�(������E��N��/�	��$
�����JÂ���X��@�nx�T�$��J��r `V�3.��kq4c��kF��tX9����W��-��6}��	�O�v�1���і�m�Bح����Ѩ<y��֮�ׄ���5��-@ai����~8Co6z���9[s�^][�w�2�+Gt���p7�	���1�ۨK�{�'RN�M��e���<4.�h+����9�A"��'Z~�ë!Ѷ���31H�/[�Q%+��h��az�)�6gH��m�z:�v����|�A_�)0�/AZ��n������M/������	� ��]�ǂ������q����R����,y��m�ӛF��g	�7.�|���y=	�\�Jc��i���˞�DZ#D�L-r[ې`��4��V�=���~��k�� yK��fڹ"��^�I �F��f�au4�Ra����C.��'�D$�w_�FT?�Z��(`�T���GS+�	�6�K��YV3�D�*<�h���v!9�\M��ǯl�0֞	�a�p�̦�b�I�BM���H�[o��Y��'�x�wr�e��(�~0��,��ֽ��:�
xr�%#�<1�K5��e��
���bW�vy&GJr��jz�[Rg�\�Q� �u_���|�����Gv{��TKwp������lgV���A�JH�Y	8��/ݖm"�<
�(x���5�ƪ=RL�pp�g�K|��Ã�*�-��^���J���$��-Pn|�W�tHn�e�#�<� D.[�ô�A7��*�qvQP����Z	(��5ڮ� �s#����܈�8�eሦgŐ2�`I��5�a��b�0�JȖ�`�n��f �f)�I��0�ޮ�+��A�a�]��F��0�g��2��*�^;�My;�
�\��l;��5r���T��9�P"S�g"&4h���ܝ?��ϏZo��(Ŭ��y�+js�ү �Z��_�P'r`�)i�����Pm���O�Z�sֽqE��*d�Ð�D�9��{���3���[v�-�{F��c���m:D`��km�N��sԗl�8�m��_	+�H��ƹ�+��L��_�����*`�T�'�I��j[�^�i���1w�"е����E�4��y��6�r�h�[�%8�7ŒdB1Ԉ[�9U��gMC0L�jHtB�|ɳ��R�Z`�Oo����d=�$>��zK�]y�����Y�2`�8FG���'�ޕ���-�B���?�吖Z
����~���׎>mi%���U��:748��CUJ�p,����MVg=�Ϫ�����R�����@�Ќ�������3(C)�~b;ă���m���=I�����vv���Z���<n
�Bi�$�:u6�������@?UV���'r��p�,T�z�K	@��	�5ڹ���Av<I��ѥ�i�*�E�"�&�*�4!H/;L�i���|��C�8�SWQ��hUu���Z�֚&���:N�n�z�A�hF����
�z�AA��ӳ_kl�{AjF¸6����p�ez�џ��K�q�bS��y������s��|L7�eZ����hnk���4/�*�%�])��(�͵ x���pPX�HhU�fmq��������䀦��dVb�p�2�y!{��=�[�6�u)�7S/:���[�}>��I yd�Kf�آ�DɓF	��g��w��sd�$<kd ڢ���M�� � �.,�,���^:��pe������>�I�\r�P�=��H���.J�U���j
=����"�/%s�z�\U�ԙ!��ۑ�˘�<ٷ�X%���G�+mz&/b�|/����P��}�[�se/H�����&�1�X#<�v��%O� �e�Sz��?%�\?ߢ���j�֓��1i��픻D�a�p;��7�T�Y�	i1��z������Ī�30� �0���v�� ��h gi_�/k�j�^4�Q�</��WZ9a���?�@S�<�5[CH(J�5��#�6�ݶH$�d�/4�H5��^�l�rD�'������a��]����D���2�!�J��듖��l�0�az��0b�&�MeW�'��y73�Ah��s���<{'�{��M$�(�5��yS��{0?;��T��yA�wn��޺X%�Y/x����=3z�|�IL�d4fS@P�#Q��XSdJ��~:�d��Z}�Μl#"!t�G����3�ͫ���f��6n��b�Fsfi��]��c_����S|SɋK�����*�ة@�ԁ�7�I�\8Cm:iP�/Pf�Z��L;�