XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������V(��w_��C�6A�|O�n�����8�ɔ����ͨC4r�F*G�)�UqyY����d�O����(���*Lj��'�>�G^#�������p%�xG�a�.��� ����}hͩ�#S�N��Ȇ�M6�|�b��ɒW��NNF;z������i�3�E���|`_��M�
�n�-��1ѩWg��)���Ch�^>�*�i�������ǣ������Z�����q��i���j��J�b��@|��Y��f�]/Yxq�pN⏔�d��1_=��X�ÈW=nيK��߅��wL��c�mH-i�|�w�Liů��m$יI%�s��.(�Ϳ�@AZ���.S��卺b���C>�l���8�V0<)0��[�vG::��*@o� �w(��;�W;��k��������cs�f͕���ԋ�9m:lH�dj{��trf�/ɚʪ���c�Wβci�Yd�۝���OOh�5���,��H�7��������>���}n���2�E#����5��T8�!��� �"Z�u/��C�Z�,"5���\鿶<i4���&��3dWZ1k,.u�{�U��s�q��h���?J\G{���c\RM�~���vVJ'R2�!I/��?β-�'ż��?>��DO�97�)�r�u;S
���i�B���.�ޡ�`��pMT_:�ͷ�����M{٪�Y/��X�UU@���k�q��RZ�ዔ��Q�]XlxVHYEB    b8a6    1ac0�|�q�!T�¸�y������<���.�}M��2� �9��uoa�'�d�t�H�@ƌ�%n���X�:
+@�_&�y���M��wT��}c��$��q�̪=�@�����TM�q�@_��7Y�������g�����m��#Y�A��l�PBM/���#�^�	�n���.aw<���ټ(�;W�� [b�H�͚��_U'#.sa"*�%>$���~����/R3u�����-R׸�Q�Bn�����.�)�-=����"�05R_�^|a*`��~5$�3�w{�^�hBI�Mbl�g�-�U��(ӰL����Z����Gcv�a�t�,�{���r,��@��f�n+c�).��fY�Y����@p3C��&(H�e�G�l<�3� D�\_H7�t����������	eɋJ.��Y��$��#�)%)�l��Jl
�/���8r1#e��I�;���Σ�LMՊfv,>��-w����5ւ
H���$QO.n0v�i�RM<O���5��#6�����A�"�-�eSZ��l��Sx'r	�����x���9��;�5�N�!�M���!�A���΃��cZU?���H;'�岟���jY�u�fIuB�?�6,�[��]��i�'rh������*9*?]�ë+�h�e�t�j�j��1s+��PU������7�^��Cl^��}+�z��{��k��m���~qA�Q����=�ƻOw�(-dG�O/�O�|��Z"������-wWM��i��n_�P�ۍ�`Ո�	5�����1�Ex!�b���4uwU�O.��&>��Эp�+��|�*���+(�kϞ�q���*�<!B\��թX��Gt��k��19'���W��g��Xr(ݿ-���U8�
 ���� �|�*x�/9���j��OlX�]g�R!R�}�tBs�Fj(��Y*���m6F�ZQM��i�|�_�x{��F''���W������Z��
^w3���MOWjx�V�5����`"x��֢���P~Dd�I.�P�+-AP�	�ˆ�s���=Ȝ��ѧB���>O�,$����-eG��<���5��Q<��J�ZW4����?�P$ -k��YR6��~�-@̟������W�� �-�ǫ������`�P'��,O�_	7�����}<-�@S�O���[�ڨ��v�����U�.km���@���+���}��-9�YPnH�O�*:;]�WS߹�����x�/�܀I��Ҽ{P���+����ƍʴ�̚�������èJ�«�^���䐸^�9�v�O�*�����&2����Z�1�eO$�����2�`S�L0C:���
`B�E���Ik˵&[�ZH���ؑQ��8�Ua���<6�����Ĝ���Tt+Ԯ+���(=��QP�����-" V�H�����;�T���d�u�ǿ����SF�S�����kDI�`Z�6� ����\�	��N-���Y�9+�N�bd�G�Na�{��y_��ª0%�����IST����Q�L(*i��:~�:&���?#��ʨ_R�-�o�ߛ/��<溔%,ilU����ʿ.�3,9F�f���P����k��W��s�28�f=��M�����^u��y���zAe%��l��<ʑ�y5����5��S�Q�����:m$]�ڊ�1�P�*��կ��u���T2h�ݣ��Nl@�5���}�8�1��l�Z�/P�xN��f��}P*�����^d��z )��xn`Y�䬵�n�.�!��͜�)g'��QN�[AB��f�]��~L8�ɁV&�kf7r�g0:b���q�Y����lh��nl� Vn��s��V�"�����0c�#�a�U��ښ�R`�m��y��o}-����[����{x�m��Hc@�8���i��$\��^���"Nۆ ?������̼��A)������$j1�qi)]׺W�Q��8U����Df��C�'�Z�%��d��Y�t��� �s�m�����������dyq�+B�eˁB�Ӑ�Hg����y��5RTLbg s���e���S�3���U���U��N�U_�w&��ɭ�,��68���&�0զ���R �2J�m�}·�߱�����H���|�#��
 ̠��_�p�$�,n�5c�ҏS����r�F���E>���>��5��q7��:�T���N���qhkPo�4���1Ɏ�K���N;���8*�K	�yW�)�>e�A���Ou0d6������ʒr�]�W�n
d-_����7xJG�%�q}P��]Q���A����'=Cd[�0���F�h~�K�G�y�����"Zm�<�4�:H:DAʂ��~�}�k�:�A����Z���D��>-�'�@�΍H"D=E	`�+|� �F�P��N1��������6�r�UR;���O^��?��}?�U����xAV�Ɵni�d�$�Z����e{3e���qL�n5x����B�B�ꔜJ]$h�4�`җ�x�X�T͇OY�k�%�$)e��9���__ݐw��"����$Q�nP�?XJ�L���
꾝Zj�����B����D��5��d	k*�.��[TC�����2{Ԓ�<$<FGEmQ��:.؏N,��=j�P�z������/N�_1��K�Y�Sя�uos���|V�e�¼�V,$��R�> <�����`��FSqBh��;�AmA���l0�,���+�%�)Mg�	�l_���O���G�Qi�׵! ZI�v��ԍF�lp�2�kת=ߛ�U.�c|[e�u� �t/6p���i!�2!"�8�0�ݣ��K��Q��O�����J���x��TNu9���{�� տ#V�#Kz}y�j���
�v��I����@���<���&��A�䯵|�m<3���<��!�K�e:+m��*W�F7���"���������"���������l�b���8b~���ʳ��� $+���S���J���q$e�qm{lgC�_�x?a
��u�k����ðխ 8D���`FB8�9�]�0T�<��ȒP
ad�l�(ޞ��l�Y��I��v�˔�J4C�	�l�vg{��k�p*�k ,4�]�p ���3�\�wXa�-V�D
#��\���!/ah:��'���g���_B�R���!��=LS b֖���F�ֳ��\q��qX���>�Z��ޠ�_�^��w�>�����78㳟}�O��/�w2x�f�:\�\�R�Q����<Oq0�
z��3��SBA�ENӖ5�:���^=h�Hx`���l�:��d��vm^	���y����oGt��;�&}���Ξ	WQW`$]�`aN�A�%h34���J�d�r���ܳH�D��'b3�Wـ�m����)a4b�o�����dp��{�l��{�>/y2��P���t����+G0�������S`�(VQ7#�lΤ�m}��찍�����6x��{# �V�v�R�H^^�gs���L��a�4pP��޸��{�KT-c�p����ܑ �̷Ŭj�؍���צ&���K��d���0�F^��@��}�7�0��]��oeY�q�������HI��J�b �}_^��;U`�3u��q4��r]���m�>ݞ�>%v.�A�Z�5�#?F�YU���%��tT�_ht��<���u�����b�J�Q�[>>��/JދL4� �����9��GW���X/���y��c�����t�rR����a����TK�px�cU*��¨Q��xU��{�.��+
��8ֽz�2u?L��¬O�n���#E7�M&�B*���0�"��q�1V�WB�}'��)��˺��CZ�'�z�9�0�K�L�3�����j@��m��̣�,���Y!',¿��qhHM[���;-�#�r��r�����`��[ҡ��?q�l28��s�cY?�FWs:S�f� �(��?k�e��;����i#:V��T�Sg�8�U+x�"��_���'0(��k������Rq���GV�ys[�V�&�dEE��$y4+_�_�ƔG����!�ɥ�l�1_CTzA�2T'����Q�,�W�7��kl�C8���F�'���Tl�Ng&�����	�J�ƹ�}��"̙����IM`M��0�*���Ffa��|��N]�6E�����d���`60�b���v�s�qka����g� O~�1��{:�@�)���D�ؐª��v�I(/�ŦJ�OZ�8&s+��l�/�j�K�L)D�j
�?����[o��OH�E���'���d�-:���aSt�$����!�
X���=ɔw�a���*<�:�U��d6I�d��^v�kA�oA�8dX��NԈ7e.'A㶱Q��7V��s{y������F���WO?>��UzQYAM'j��G܆���7�7���)��]�P���_͞�����Mi'�è�]�Y2�S�w�����6E��W:Wx�֪�DO��=�=t�
=N>�VÛs|~I���|*<��_袲�,�ۅ���� n2p�t&s4�1ĝl�'GQ.H�gM�7�ΰu`���"��[8Bā�a?�oyN.`6�uh��`U�٥�/�y�_����&z75o���7e�C�Q��ch�L�5O�^�
 <�,Ĺe�GqN�ox|�ȷ+��o�w\��� t�O��5���+>�GoVZ|e\f���zo��6��Yֿ���!�����Rl�n�^^�iE�ſ��k�A8\�x}!� �廫��̓
G[�c����n�������ܚo���t�' �� ��=M�;�Fu�,CN��!�^�숹����x,RR&6d�|"0?���cHs�FB9�y�g���K�J;,ҁ]:�	��E{w>��+�@�I#��"#�C-B.�m��^vϔ�6V]�Yi���W��E����Ah��������J�������+�)�b�z��Kf�W��HB�!��7����*\*k)G<湐�+Bv�L�}�_�ӫ�*+�)`-I�(ޛ�[}P���������:ߕ�v�G���`�>o��u?��φ�
F�X���ЁtPD�+�92�#x{gDҭ�.�-��<�n\���S�p��D�����mف����&��,�׳���^^涹.	ṹ�Q^��Ҙ9��ۀ$4 !Z}��!�$��fm�Y����Knڊ����'�t��m����9���	�>��I���]-M\�p�yӨ��C$89�`�i�1(�o��s��(�{�	���A�|��3��I���pb(��{�}�?��s�5�B�����9�8Kk�=���wֱ�2k�HB���O>� �ݗ�s�Le8����U)�4�7+j��ǶC�0��`�	�h�@�Nst2��\-�'���̻��A9������y����8��/���������*��?S�˻Tx.!7�uؑ�擛n�6u-`��5�H	i|�ت9WYԻ[�e�r�\�x�u�<���M��T�X�`�����V	&�д��خ���X+��]^��$T����z�z2dM}L˺���u>�Uu�GP[�K�8��ݐ=�e4�1t����I	3}�$*<�Q���-x�3Y���,��E��G�C�iQD�K� �4
��:���j5�bҳZ��ța�)�.[�Ӈ�{��?��Or���+�lk�� ��ޱ�mS푺Sl��	��~���f�X�~�R�mL�b�Sh���nV�0�`��u�y}D�W.��d�KH ��!2n=!�bא�%l���3嵻�8��]�,��c�MJ�搙K�D\da������wx���GEC�,Kpk�u��w�7]'�#�k��'�H�|���s��)H9�ڱ���[�n�,0�/�4��v<+�|F�h�@%�|�ўF�/������1K��<��6޲i"+�^e�����/�_Q�."�h���M������~�?tO�t��ѐ��b���|��"њ����d�)#v稵:� S�?�������yl�x����|-Id�!��lY����\g��*.��Wv)S��M�:F�ZZ�5�=�7:N?�+��ܹ�-A�l�=��%�£�������.WUZk�suګ��n��+�XFB
���l�Wȧ�����H"���k�eK�dlPV��~��d�
�w��������ī��jUͤ�Y�E��E��)�F�K�Eߗ/v�#�;��_A� Ê�S��P�yl�g'�^��Dkb}1폑�0�?
(	��4w��9j���Ce\�/�ܲq0H��1�J�8�
+(>\C�W�?g�f"�u�0^�8C"�V�Þ�)�)�܈�OO9�ѳ �5��?PA?�p��VI�8vd���*��r���(�-�4� pv[��م�:�ފ�rt8��/��/<�N��Գ#.h3_����YX��)Z��{$Ͼ+-3�1+y�a1�	��*�۰o7�l1nʧ���OB,P"h1O�a�`�g��A���J��:��L͠����:�?ͦ`�[���]Q9j"<1�~�D|�N���m��
��\hv�E����
��='�B7�eK�@���r�8c)�M,���VR�e�i�K�Y6�Z~����ǱX���v��I�o�*�?�Y���낍�!�I�+��[�#s��N�9d*�I�5���~�/�!5K�h�aN8���V�^��c�����M�#�/@�)���_vX�z�X$&	���S� ��Gy����CN