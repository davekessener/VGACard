XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&��m�G	V�{�o�W6{I�� Fp��UV��^?���`� h������H?�B�{�~��g��n�[WR:��A����TH*(�u������6Q�'��{,�p���/��
�S��8���5g����X�����b�Zb52ȓ���&�,�N�?7eҵ�E�L�Һ��U�;縀���u�n���*K��5<��1�+������Tq�/-�F �r������g�|�~d�%�ձ��2C��T*��.W?~��{�c���,�q�@�bJcT\� ��t%���P����m$�;�
�k $u4R�����Eps]y��� �)W��Qk�Z��
+W.γä�RA 1��䷢�
��Sw�-�,;�m�v�ћ��<�s�"�`��
��OQ/)�ƧT�+�G��wetfa)��L����f�mM�r�5�dꢖ S�|0+/�L�s��jՌ��� ʋ�㲟cE
/�;=2�t�Eem����BW��l�4���v����t��n�Oj�M�#��?����?~���A|���g��/�>��7J-7���G䌃��v)�����:��(.z�)�]�8��H��\y�fQ=��D/�;�K�����2��GI�T������g .]~ƏGqM��%l��eL_@xZ2b;u	DLչ��}�C-�sR�$�d7�<��^js�0֚�_J)f=��`C��?@\�j3��|rU���jK��p�b�1��veshz۳F�Q!�w��XlxVHYEB    c3e8    1d20���`���P6=�%�"qX���5�P��e����6?L@,�zO�l�]|�^�ɜ/�ޛh��@[@Gs�'K8�V�?����|Z�m_ :�Un�@��}sO�3����?�y��1�R��	��
�)-�0Gi������C���Q��2`L��M�����gf"�����7��^a�%�j�G�����{!�A�c� t��D7x�8ɏF���6Le �Js��𱒫Y���s��,�1h�'��&���9`!��R�Q�CV�M>�2E�Z��|8�饣��E����
�y·	�i�TFM:���˟<��>�;���%'��L���o�����{ f�s\�40��u��ܠ�OiUVf��1��F�n�m�yŚSL�ʖ�W��M;ߎ�F��҄`�S��b���훽�N�;�Q:?��/]�1*0�ߠ�&��!&O ��]��[�D ��vw�X�.*�l�,^w"��4Y����^٫�C����,�@��n��� �5ZZt��.�sR�����v�]UK�42�b[�?��'���n��DU�*oupa8y�uOI��<��S��P�P�\�J�6���G�J#�� �S%�Ϝ�:z,Qt����yT��]�Z�i)e��$�p�xP&[[Ho�W�gό�a�����ݤ��ۋE2�2;,1ݛS��τ -�"��;�߁�Rz�q/RS��|a�V4`��X�h͂���k�E���s��de�����S8�XC/k=�L��
� ���fc󡖕ڑ?eU.��}�F�."~�Ot�����d�Z�c��Pl���r�Ú���S�4u�n��L��S��Ǳ��oA�c6��]�N��Pe�&=����vN5:>x���|�`$v4��S��(��	�|()��O��oR�".������zI��d�ny��H ��eu^�6�ׁ���A�Q
���2V͔2�b�A|�G�oiy9�d�/�;I'��3��Ȕ�NC��M��1h�h�kw�@�*I����׽gt#cF��P�(��UoDqP/����5����!6�r���u=��
:�.�6&�n2B�[�,#m\�Y\��3NΒ�f%�'TJs�
�e�
��H�6/��t"��=P~��"�D����y�!�]�T�T[1TYR
34��_G�w�P+h#`)i�k֋�)�������Ϭt�O��+�����󻤡���zi��*ʀ������-�PB�րT�X҅��1/LRg�(��N\	�xx};o%|ln��K�4{�~�J>Ѵi�4��z���ùk�]��������M�s�BW�&/�L��c��5hߍ�G6�6�2�3��D֐N��Ò�2���7g���_�3K4"�n�V�C~���h�n斾��`~�77��Ԩ7��f1�;~+mY��^I�	����Dh
{��27OǆK�Up;5��^o��i*w�E����\���(��s�Ds��
~�vÌS���#���GȤ͋
!9�� /y�| �K�<�w�i�!ƨ@m�����?^	�W܆��4�,� ~k�mu����G��7W�j�:w�ks������C<��z�{� ?+�mQqG���q>�z&�e>���5�tZ<f�x�#j<譱DIJ���6{�uM�I��V�U�0�lX�W�M��A���f+�g{�]K�6������NR�՟!JxH����ʵ�8"N����&i��Q���p���Y?Q��	��L��Q�׼���,������z@:����<'K�T*�ג����jI�4~0��U�Sw�lո��0s��M��e�<e�P�͉5'ey�6�N�Nĵ�����9CD��j$��#i��\l������S@^��D,qm��n�O ����a�|ӣ��4ٓr��9%��f����l	�
^�>�^���V-:�����Vx5�&x�*O��9Ϭ����r�sXX/�;������	��s��C镩|�ؾ��#�gX�����'������`�Ο`:�c
��f!ٷ��9�v@a��\FU��Nq���Kp���� �uc�������	˞����.�ƭ�����<Ԭ]ֈ@�u[����	ɋ M�I�e��v����(���ݒ�"��*ZC-r�i�
~+��9JeMm���oJ��|�T�ǇK��d�c�N~P��4e't�[>i}-�@8����	�:D��(V}Ʃ"d=��鑶�_�欃74E�#_:��$W)q8��S��cv`��g~|�SQ`�[�(@�(�,{�X�t��^a�_�Zv�ԭ�z=`4�X'}�V��3sg�l�ŗ[s[�1�o_�KԊ�X�<�b���8�\f�EUپ��Rg���I�.ܫ�6�_}i׍�.o�,�R��_5�y�(���q>�k���&ì�?9���ON�u)h��W�?� ��e�n�@ �^���-�V�8���:�(f�eH�x}����;�}�3�;y�|���>��F��
�5UF�T\��:-f=ʔh$<�}���3��E���g��t�c(,>:|��X?�ok^
o�xf~k�M9uƇ�8�؏PVI�dE8�ܐ�|��r��Ks��'hS�L惤�CKaT#N�Av\��*�K֩皾1���X����m倃�K��nl$;;7o��Ν�+���(r�W�3�D��`5?)eؠ̻F��~����L�X��x�*�1��b�X���!9�b���ξqi�+�����3��	!x���ޑ�������N^⛠��A[L�.��p:jD��@�rC��);-�3e��r���!)��o'esh~{�m$wa�wٴ�n���EK���vJW�g�7���aC�j�����l�*�~�1�˘����@�Z=V��$�|B������ꡛ2��_�7��lF�֜��a��i;��/G���SR#²`m��X���;�ŀ�#m��^
5\�jWң�)lG����麴I��"`I�ȩ��;f��̮;Kq���|�g���s����^ύX��+EL7�v�����H7��Ov잊�����-]c�CV�M�Oq����i
>Ŋ����\��6iA����3l�FcP]2��tB�CY��uYِ� 5
�*a��0�L*��ӈ����(�;���A��>k��K�WC	�ӟ���S�"(�6������^<䏱D�rS@p�F|���$�|��x�uc���/�	�Ev:u}��]DX�.А����:��TA�ZA���D1��!�,�<:=Y����F�}�A�����T���!�1�"13,�3f���	lP�Cr	1�G��f�:@�������Y�q��N�@��f�NL�_\�v� E/��F0����~�y��k+�B~OEO��b[��5����D4Ć{ٶ�Fy��q�T�����W-=>( ޙ��ځ>���ڴh1{쵑+�j�˯��lޞX�]���~�!?�"|�m��_�9e�Ve����6�<�l��8m�R8�6,x��ѳI!q�`��ӧ��>�%���Tr�M�p��aȨ	�_���>�Q��IDH�.X�̷�+�˚^���N�� ��^�?|!a��I��ud���ƕ}�����E�L/Ƙ�q(��v��b���n���B�ެ�Jq&+�k��Te�42��<2 �b"嶚�D�H���nS�n}�

�*�i����pNeIc�|��k����n8�$�K����(c-Ó&����<1�!���o�~J���0գ�`�T�k�,�`��L�P���^
W�`�\��}F1���lIo<ZtcH2�r=�G�o���w	�����\�l����Wn�N'sl/�qn�i���2����?��ĥ=�wD�S �f�  
��$,Q���#��E����9f���i?��e\v�)�C����f���,�;�'*1��֣�R-��>��m��u��ͥB���ܸ>O��1X��˚��$����_�/KW����:�5S�X��kR[yP�3�^��t��9�v�W-|���8�U�6�����y����Jb�Z�����x�3E�,��`p2H��}�+�HZ9�:Sf%�l����er��kF�����9��*/=������W��
��F���I��ig磉Ձ� �q���E�G^����ސn���p�d��0���m3���l]��(΂�����N�H�����֊�cR�rލtK���<&e����z!L��������Q�R�G��c�]�٭�s>*��6���8fp5��r��(z-#�Ѻ�(��e�Rkn���̐� #�/Ln�3�����C�-J�-�>!��;��Q�����-��٢�X�����쬴k"7�O_���w�������7��ӐX���v;�m����e���������Mq>��h��i�m��n�UX{�c�'i��j���=��:y"rܐ�w�8%����С}�s��d�@�	��O��ѓ�6o�6� �wY��rݪ�}>��z�\ �ab�
��/N��/jɊd[�FNjs�����+ٺ|R%Ps�`�	�
p�����Up3�n�b^3U�L���M�lS��{���l#��C&ϱOh�ߓXkdغ���^+f���Lb$9��/�.�l���8N�"�y��m$�*$�T�0�v�{E �O∋Ax����M�jK�NnBe��HOv��F-��ͦ>�/:�㪧�[���9с���9K��P���>����HZ#�O�[��#G�XL�9"��DR��pv3��s���^�t���B��g̦�*mk��d�kpfp�2��W�b��21{�����q%�`���_���b%�K��XA�� H�=��JXyW*%��5P��%����i�M�F�ٹ��B��<6E|����)���kR��+C�)'��f���S<s��=�vd�)s�5�f����a�0s] �E�z�2:d�/�l+�n𼡒��2�0[J���7c���ć��*
� �`����_�ț㪭�ø��F�`�]�.B�<��*�{��?Bw.�	���{:-��ep�W�i[]�A��]�_����Iu�UjD�C|��ʝ�&v:�kv����;i��j�x-'�:��ܪ��U��C�"US�HHJ+9��.���"9v9�׻b����;v +�>� 5�ֶ�J�X[��I��Ny9F#�>�W�A�h��t5��������oOц��.0.�
���{��p�E���t="t �k�ǯ2 �X
�]��{R�VL����9��k�U� ��8�I�qT��p'I�@d�Y�	� ^����U�g)~q��X���$�����d_3%k! �	��Z��Մ�wvel旴%��s��e�I�˻��'�e&0�7�!^��V���V�ԃ-v'���f�M���հ���h���#�[�����B�[N�	#j=#ɻ�+��y�yü����ٹ���$������l��3��d����yO ��Ȑ"U�y���� ���Q<e�1z�{�
E~co��"̄�?)`�
Lw���o�hю7�H-�i���)i4��K�P�w��F�d�9Z!IT����B�W�h|;ay��y����\�M����.���Q�ū��H����:�Sp���ό��e��� �Q�F
����Z5�X��?l�!�s�����m�E��r�,D<���ȑ�H^��f���"W/.<l��ا�M8tǭ��JIQuM�_7	��{ׅ]Z�Ɉ2��8���;r�c�q��=��Y�%��4�n��Ʀ�L�י���LcX����h�3���������E1&A_��<�Q�T���F�-Խ0+E
P�ڠ?i�>��75�ŠE�Be1�	��W��9&gU�Q!Y l������oЄ�"�tZ�iC��5 �3C5�rӪ��T�̣��j�� 7�5���\��j8�E�O��~K��;\��8�}#���y0���&l!����>���D�/b��9��yx��z�B�k;ۋuc��	��`�)P�+�B��?B�첋��OA������m?FKe^��F�%������C_��4$ίǹv�zB%0:������ɶ�8�}Q,^)���o���I�"�|���䯦d\�&�;��qp��*������s�_I+@;���@�'Y#e��OD���rAXo�\-�/��mf���S�P|��ŉ��t}rc��`ofW�����:=�h6�Ӈ�iK֔x��(xT�h�畼韜�N(6%����F�5���=[kz���m]I,t�"�l��m=�V8F�|��w�� -`dkc���72r־��.ф ��u�e�V�ٌ�8��Y��=�⁥�iz�?|����s�m�.���>�/N9��a���ɽ���i7�p3V���9y8��f�Ǫ]it�ϧ63i�-�I#���؀l���CNk)l	8���-t&k�>o<|��t����h�ڛ<N
4M��4`�| t&�s�Ns���i��1�� �N:��+S��@Z���幞I���u����x@lsKa�#�����ů�YS�,S��,%PU�G�r#'���/6�:J��3��tɼ��
`��c��S�~��ak���X6ۯ�H�|�+7	հ�����S���a��"L���1�)�N]�UE�0�u�:1p���gs�ݕ!(]x�YP�XI�]M��`�D���X/ą�;�ґ�&�����(�+�6)��Xh���:�BJVJ�_m��ۥ���s�q
s3v7�m:g[��e�s��,,�}�u�`|����qk�䆶��n���9�
��o��A߂1�&�lL�k^F9�e���U��8AE��GR�z-�`�ˣ�,@c-���5�o���k@���t4��S]����e���W]$�n��l�{�G���<{o���s�Ԩ//��&��4�a*R�(g|���17��4x����'�{�HGdnۑ!�[����
M{����{^wFG���ǒs�/�Dz!���n��p��Ե1��t��9!0��Ԋ�*!����\7�*��.x]�Z�OŨʶom��ؓ��N�[TM�f��5u�=;b����58�%J���9%ɧS�;1A�$U杜�;���9��?�_H��:��1� �mf)�IY�V�m%��)���xTa3�3��I#v��d�|4���[j��=4�Z�����/ �ƞ��"�/��Nb��*��&\"���fm�mhdҞ�3i���6���e��	w�	
�c:��W�V��)WLwı��e��0/�j�4�Jk#��lz��L=���A������0�1��L�]W�]N҈�L���Q�7\.9�g	>����?2iY��?7s