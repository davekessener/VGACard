XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E(�t0��֠���8ZQ�	��V�X�`�2i�����9��R����T=n����p�� ���Li�=�b�{��LR�V�*����!��f!��~|B0'�z,��iW�)TL�m����5DEۚ��e�O*���V ��K�9 ��a�Adg���((+�P��>�aM"���D�U�n�͊C�t�!��i�*y�
F�Y�-�
����4�<��}pI�B��~5�^��E�A�AuN�=��O����k��\�͠��=�y��C��u�`����Ύ<���!R������~{N���T��uJ(�?)>(ot��²��. y�/�S����T[;��a<3G�t���U�z<s��SAO(�[����,�A��kI�}����4���q���\KY��-ÖɃJ=�:�e������/1�ߎ���3Cjՙ��֒�GF�y{wL�:�0��r��`�v�b��;�������ud���pn&�$�Em늓tL�r�G >�^����cS�pJg�1,��Gd=/�2�ys��	ܕ�S���N�C^I�*<��,'��*�\C�v+*y�Ow���.]�p�;�O61���fO��n��
4��gZ��1�q��K?���jd7�&=t8T��H(�@�S�v��z�s&f�]���[�d���.a5���0~�dﴇ��z'u����#�l�)zx֚�՞D<#j�_��/��@[��F�@�Tt91��bI�/l�&�\'	*u�h�Y��)ZIRBXlxVHYEB    fa00    2020'�pbFPz�#��n�"������_M�}���"6�n�r�Ob�ۙ��U�j/�ê�u�}�`�T���\��u|��;��tyGoԹ9����y�y�i�we/�D���e!R���|t,C�� ��nh8��K r�~^��>߻��˘�'q�O��tE)�$J��o��m�k~4c���%���G�/v�$߀�����:h����`��,8�D�Y[-�YeDc�������Hpm�afF�jʥ1dB���,�~��:䳏��9h�_I�%��J�M$������EWm�9��h����:L��pb�YI�����G\a�o�G�0�@e�[x~�DF��ޯ��.����w��m1r�ܽ��c[��/�z�Bs�;rs����*��6VoY'2BV#N�B�������: �6ﰂ�p��BзJlx�=�,U�h��tqU�dhC�"d�˃HzN�p���L�pd���R�v�Eow�ϩ��W7h�y�f�O�q�m�AC��3-tZgP��8��KK9�eC�]FDE{3���� 5����:z�JȄ�:Fd������&y�l�󘆖����2���)�#~~cN����C�b��/���Baxr�y��}2U5�N�l%�5q���W&���bh��{�["�;�|L�����fmR���_s�k.���M����������t��CLy?�q�T#[�4�.���I>���r˺�7PSҲ��Z8|65��.����ˉ�4D�펇5T�w��F"w������+�_��M7�K�o���"< �g�P`�|I�̻(�=<�O�ױ��0���l� c u�V�{����S�z���v�֑�h�i�G[e�gc�
fʗ��9L�({�k�����}�x[�e�`��ɽ�1�J�ǯ�5}|fQ � ���x)VJ���f8�4,#�Q���}�[�:oJΊ$��U}	W��W1�R8�?uf����3�=$ł1�-5�*��$K����ʐ����Ԛ	�aj��8�W�}�R}u�7Y�Գ|��X{��m$)��W�� I
]�~e�>�#��xu;���+����
pw�J��X�J��@�̤W�6�V�g���C�k�I����]e���a�T١f������?���,���X&i�p����$Q@"�O�&��_��lWzI��*�f���lnY��rJ��m��L侮S?�L����5�.8ݱBllf�g�[��稽���'��6�~���W�������}ɼIOj��2F�󡒭� ����D�̥���R=�A�2 �?�KWɮ��X0W#�'� �&j�]�T|F�V*�2p��K/& J��X�ZI�zy<w��V�߀��Ζ���F����~;3���K�2ޣ�*f��H����o����G1�6�V�W	����J��r��F����lL��1�#��?�ԋ�Q�Sa�U]�)y�,!�&7����]JM�]��8,�kěT���|%i�w6��i��[k ��L0��j���v�ۼ�	�fk�L���[�2�k:(W+�@������.�j%3��c�.n���d�vW���~xn��l{s��B}�0(��!\�Q"���R4j�Fe�������#��9���Uw?���!S�k,�&�F��5X��U�����z%�/�e�d*G(q�7��8����m�杯K�!ZTܚ����xᕢ#�G�3��+�@��y��8r��uNk>~�r���9�t
zɂ��E��&D�NZ�gi���\�)~u�B����Ix��3Y����[▓|O�@g��J����˼�44��zz����^n�k5Y���7�ɯ���b��R��������v_/ZRy�v��V��+"X���E�G���]SYt��$p�削��\=��C7S�7��.g)���BA�m��95B�/�����)�ʁD�b"��w@�si��S�����cǫӅsl2���9h6��f��@Nϧ)�'I*Cw��P>U��7��e*��@�R��n���6N�XGƸ��K�U��;+��\�O�hP�t�[<�(=��0c�ڸ%�R����Yr�l�=Hp����:�g08�{�C㔳"�n"{HA�Yg�ڨg�����|�о(ȶmn)X��7ɐ�ka����h�o�����8֧��&����<��FkZEpC,Q�$�:+EF%+��Vx�{��&ׂ�O�a�����A�C��
m�� ��y1�j,`�,��[*~��Jk����:Rҙ��4 gA����׻�e7v�F�-w�7����&�,ن�*jh!Z�p���{fԅ�f�w��=,^��
�\�:����^���/�l�	ґKX^j��(ĈG�|�H�~�v�TD=)ݤ⭾f!V�x�1�i0z2��ZǄM���}�l�Y�*~u�+-���W�/#�`�� 3��Kj��,|�Y�=����R�R�
��[�_WD��h;�M�)x{��`�ų eH�����5���]���KW���	j�>�o�}�MM\ī�1Gh�8��B�3I2M^Xr�"�/����8�����9I��FYW�Ī�)E��qy���F\�Ua�+��қ�����A��`B��Z>?7���.�_���E�n��0�|��=4Zɰ�J( �H���$.�N��G�nG���|�;��(�:*����<�91,�;��(���<��Z;���A����v��Z��m4EX�k?�<h����:SNA<`
��\% �Z��� ��Q�p� ��~���+�6�@�\s�����9�A[��RB(�tk���ܔl�B1�Sv�.�t�W���:~��׹��Ij�GsX���(��pT��4%��I��rpssb+!+�h�%��R{Ê�2�|돒�zΟЉ0r�pX��i�i��7��<_�-d�h���s BBr�U6�����Q�ef���c��I���A���4��؆
p�U��#����zB�ODg[�c��)�o�V��Mt�gH=V!l��)~+zM?0��e���x%�%�f3AȽt��⫷,z��ŀ�+�ʘ=&�5�A�X|�Z�&�Co�'e�
�(@#�[ ��D��Ap�%r��9�K�g)	�����z�����V����>j(0��e|rw�:P�PIL�$���p� ��\�Ew�璘�%&xoWtLvp����r�g�ᏌY|���f�y��6x�7�{�'����2w�럛GIS�ZTyb��.r}�<}����� w�bh�4gAѼ>�	X������T_��%Ц�ޕ�p�c��p�G�c@�e�zDv>���ަ�p���֒f�FV#�9LfV�e���������S����Z*�C4+��ū�Q)G�A ��C'Z��Ĩeh�8���X���|�5���i��]�uWM��cL4�Th�Q;ɬ���`���j�����E1�iz����` ��l���/�v���}q��˾n��c/�']�v��ŲS��s�>1bu��0�8�Ѥ�
�C2��z��Ů�����ԎgS��u@[?���F�LJ5�ܭ0�g�2�1>��)p�-R>��[�ܒ�*3�K$�5�Y�)�ŵ��ѵv���t�d�sd@������Y��4-�E-�n �9�Q6	 �뢀�Rɜ�^2��Z�Qz]x���l��q���Ù+�˯@��lѳ�����PH�4�$�J@��^{} �NF`�s�1�En�פֿ�+�JJI7q�;~�)�6N�Rf;�:��d �	~�ЂA�l"zevJ����L(B�M*)*�7�։b�e�	��^O�����=��̐m�L5�O~h<�@�t��Us�ѧks*�x��a��A��!ז�L�����=��FU�ہ����0q��oK�%��l$���k����l��T��2pC�}Q@$1����hm�CO	�3��C�! �Q�gO?jU�Hj�p�Y���7}�d[�s�*�{'C �+am�bΎ�q�ʫ43c�~T$����m��~�D��q%pU+��V����WˈP7��v{���*�W5��Q�u��Kk�m��ݧ��0�R��ڮ.��na%U�ְ�b��N���D��2�ݶES'&����ߝ՟jԊP��I��B�+��ZQ���޲h�є�A��{ljI���-pS���I���ȝ�ٓ��5��Ȥ�\lv��~h��ڢ��C97AʱOyi����`��"�)fw�(�ۄ�%©��������UJ�Y��c3�a!�ʠN���>x�JO|C�,��Q�����۞8�
����`y%����^�Ve��-�M� 	k�|��gT���ݠ���1���'m}�B���"��򛶒�4�W{��l�p����}����fil�RQ���-oGWǼ��]9���8��6�.���?<����쑉���K�{������{��G�ne���4Ѷ�X���.#��B�K�K���L�WI�LS�O��ɍ���`�r����Z�a�p����x�!ꄝ�J�
��� z��[�x���|�GaD���+�ݧB�vw>����>�x��p�Z��BJ�(��|�ϭ�����l�i���I[1����e������f6�����L7��M�����.���1{�zwZ$�=��A[�B�_����GY�TȂ�v�q� ��z����E~��q���2f���
d�e_,}�x�gA�&~L;�6����ZQ@��t[[�LRow&؄�)4�K��FE���ƞj&���:�j�����e�>��0�,�g�p�����+��!0UU`h�W�	�0j9��*9��
����u�Ї|���+"u�g�ݝ��+qQ�$���
���V�J�j��瘈�����S�PiX`�]�`���[5g�E)Z ę��۵���Pa�Ȣ�;|�3t ��ۗPƠNo��<eM���>�vM��ڦ <����,!������ga�<B��$G�ȥ�mƺ�ٺR�V���aD��������~E`,jI	>��)ϟ�K�9�$���a^�.��W��:��1�Y��N(z�h�>]�ܨ=�m/����i��8)���Ҩگ���0-[�6�"�%�֊C1W6���j���Ar�vOq ���H��-*:t�q�M��:S���7���_P�zghhg�cWT������w�2Xz��5�U�<�uX8��Ս��M��>*�4��X�üES����S��BJA�ԍm!�i��	uP���9�[[��ضv���6it<���ÜW�%���%��K��M��u�!D�w6�U�̙� VeG5�cS��^:�sg���j�ڙ<=���:7��K,�W��ȥ���o�m�0��-���.���@����TIy��C%�^(�.nI���J�ov�ļ�4�Tʆ��o�.��f�M���s-��v�o�;�0��|C��%� �
�;��t���ClG��R�N˩���i����#�$�B�'���aRoQ�j d�S��F�3�l})R�I7f�r!�|}��
<϶�~�f���1��K����<�;�w���W�	O�5�Q`3�k�;H"�u�.D��ۣ�L_����@:�h>�Ό��?�t��Hf��q�K�D��r�#&{ސea����^uIW����u�r����S�h*��^W�S�E�۶jɲ��	�*;S�*������k����OJ�EN�;ҰS��^��O��0:��m��͠��D9�K�,ur�e>p��Q�ٔ���60Ş�$�k��!;����n絻�a.M8���)�'&� ��z|I4[j�}���p��B3v;?�ʛ���7a���!��38)pF��.�ɫ�͐�5-;�B�	CO���.�������E�kړ�b�.�&����m�$�ݏ�V��𳖔/�M"fK�7*3h�­q,	K���^*���1��̺��d��,KO����`b���:P�c�O.yH�S�<�Z���FZ��s��Aȋ��1�*�ë�1�jɻ���Д��<pQd�U̱���ԅC!혨�����ZƓ;!k��DB�q��Xj��ѵ*Tg�慉n��B3���K��t��Y��H2��f�؝S\uT)��#.R����5F��1��q5��<��B���<C{�-r�C���/S�ړ��Ny�V���ݪ
��,fv�t��	w6Ց��"j�c�`'/Ju��M�R��p��e�f�PJdW�a�ˀ\V��G1����).��W��=*��L1?.��9�+�����Lأ��^�b6�?)��)\ ��ibK�����s���L���<Ke�'`s8�}%�`�wI�������6�8,l��؎�\F`^w�}�w%���p���9�. �אS=鎮L���x�
��T�t��w�S�@1'�}~��~geDfJD�p%�ޡo5@�d�=����L��=���6B�=<���� �4}�q�/�[B�2'8k��;5��0u���Zi�Z�0��Į7v�,̼!ډ��"���_�Z�A�`2z%��*�.0��ߒ8�󔯙�KL�>^�����D�A
{3�K�q�w�����e��ƪo/�����d���� Mj���_�D�1�X(Z�Xw3� �k{z&����X�M�,,�X0�i���^Nv/!v(@i��3u1���1�{TR�������RU�ǀզ�$7璜��ݪ�p����A��A�6莝���G�3X'�KFFuUQ�E�s�hTBv(�>�`<֭U��88!<�rl����F!|X~�ᩉų|��.�200g"&�/X.\@r����/]�dP[��3�yNzz�q��vυ�U�,�E���l��k���\��}	����v����H�^�p&�L�m�!h=��ߐh��D�ZE�&�����]-��[2aO�_9���77�����N�q-�	��Rt[�;�N�X�2��	�i��x���{9�>�����`�KV�i��,� �"� ����Qr͜h�b���ǌ�b[��.`e���>���
���SM�g������կِ�Uݏ�	
�)��sVaK�]r~�j?��>:%��%�x�vu���m��o4'Oٰ[ɏ�	��F���Bf<CD�N�#��0�v������UG;�����EYe|�@lB�+���B�,�����X�y�N"J�=d��Ι�>�A��t-�)���~~�/�P(�:-��?�P�����s� m�7�&���g����� !gӎ�ً����N��uZE���3CҞ�輷;Ƈ�iX�8+o�2�kY>�n�x�2=�� 9_?w��QJ��Bԍ��Ɂi sjZ}�D��L���W�3+�P������{�I�����Tem�W;�+�Q5xz9���u��f�3�$��E7����`P9@��K[���\OPWV�ޟI�/1�A�(��v$��=�:2I.E��ѧ9S��йN�g�]=O��Q Qj1��&���\�\��/��LpJ�҇���@߫�T����0e�j�'x�J8����Q�'}�b	,�6��� <��
�X��Mp8�;Q�����	�1X.KXl�u}&M���x/���jAo|���Kr��K����8���;���+�Ԙ4?��_`V���[����?��Ȼ:#�ؕ""+Jߢ��q�5�Ͳ��<���@���h�>���>���;�����`���A��3|Bw�Cs��=���ma���E�\���l!0�N�߈�,����{����]�ӯ��锫�F�6���S��T�j�+�7��ch�k�m�q�ژ���eC9i�w��?�h���:�ƶ�%�\ȯ6�y�Y�?&"L�C0��-C�w����ЪHR�ۨ��e:�3�M����䁘�Q���Y7'� ��c�x���y�C�kxԯyw
���t�bM���	���oBt�w|�(O�b� �֓]'��l»��2��E��
�oIG��q�%�� P0Nn/�͋��o��ia&��}�u��#]�%S�y�;K���sK��0ڈ����e��B$��~s��^���u�^�ݤh�;ɧ���v�p̌��X�z��Ǒ���,�5����N0��H�v'���'R�/!̰�&	Z ��y4BY9��O�/��ʢ&l����T��6�1���ߤ�'�@e]�Gh�J&Q#��1�x�XlxVHYEB    cb82    12b0��3
Y",��:@����#���L�E=�uxO�^ J��"�Y�1����7귔Z\���JMDmCWw�d�HG����� ��6Es��1mE�$Onނj*��jm��
듊��25�冭��+/q��������d��'�ެEо��	�%:��"H�U��aٹq9<u��X8��3�2+�,�LQ
�������HY�6�략�p��	JD����|@p��}u�9W\�tE�C�j������nT-�D��)�V�{��.��,\��I������+����v���A�j�j��*:P�YߙA�oT����H[]9�^=�w�`�ps-��$�|	
Z胸D�]�@Uܤ�K?a��纣�	��bc8��aA����#dK�(�4i����̻����,�Җ2�|�6���ǥzEmT,��޼w �+_|XBv��n��D���,1I���뚯jr��Js��4��iL�S��GR��e��_BT>��ݖ������|�%�LJf�T��׺|���1�Ub�Q�_lP�Ta[�vR�ʉ�o��U�g�In��0��"9m·��Z<�3���r�*���]eSV_k��7���=����\a��n���S�=�E�>�i����^6R�xvQ*��������E/�i�bw�����8�ˢ��!��g_�n�g����ԕ*�G?L>� �t���hs����b�]��rK���m/������Ө@o@�~����Hm7V�|��fӡ4
Yd�X3�+K�l�z)��t �#L��鰔�}�eZ<���W3��uSp]�n�[A2�*���}/J�͌9��e���s$/�6ѕ|�6
ɌP_a|z�VK�B�z�a��K=w���z���z��M�'���D8ͮ(�&��'eԒR�;�J�xߍ�����>�Gm؜�o�U���f�=}n�Ɔ+�|F4�u�&��E�H�0t�5�b��M�C^�N����-N�q�Ky5Д��`9wq�u�+F>wKY��M
Eu��<�:h��	.S�Io�:�����R�	H�ۦ��򡨋dV£���\��pD#��|؞N���z-/�l��U�Q6�O�W�um }	�M����Ty\&�!U�4~�,8'3nV�]��>����Ք����䏘7���2���0�r.�������6rod�5�6<�&D����r��Β�byh
_�j|�-T�`�_`F�83$������+�����ut���g���q��j�
�KZ�}^7zI�G������I�8�׳�����FavY�	X 	����0�����Ni��8*4쭪?�e�(|I~1}v�~#^B4����17�:2\ވ����ֳ`b��cPP�Jέ��)'�K�i.MK �8v�+?k]	��W�b�ʉi.��5t�t�@~�)8�5h���)U"�ƮO�g�Wh�p��d�f�":��|����p��/.����-{{2M}'��Ф��p�g���=OZ�~���N�nc`opf����I�_(����;����u�$%şK��~��_��/�z�����k���0P>�uN�=��O��C�%�/�Sb<�P���R$r��/�
AX𫸉d?L��j`py�E#`�.�&���<Y�&�y���Â.1\��ʍk�"p�Ab���K���g�Zo�/Sp�ě���jT�Ϗ]��F���j�;:fY�#������Rl�7�>�i��� ��g�����O\�Zt��L�G�3[:���}�8C+�c�2���+�����k�j��=�e��~�a;I�GP�X�����qu"����@�w�.�2��س���aQ*��6�*{d����n��Wj+�=yt��76����	��)�ױ�@�
!�n.U�2��(�S��Sp��֍��ŐY�y�0�'�s6�M����o�����_�?�n� 2(h\�)�ɜC�����6�X]ęt�����θ��
�CK�~*7���I�Cb	�d�UZ�-es&Y�O�*R�<=����>�0��L�-��0N�6�F�Y��r�}�}��X�N(���䡙�m�+#�D�V�� ����$�$j���Po��4��M1�3����Ð�t>�;���}�P�{���L,�
�E�����tـ+��>j��m��2�R�K��l8� a�����.����[��{��z�kd�TrK5�X�@n2E�QY1	�b#����?<�N�F���t�)-�<�<�i2j���af�x�@HdÙ.��7�	Ka�ֺQg �����*�O`���?�IG�ļfu���Il�C���b�\h'�������v�����6 ��a!hKE�T��p������
�٘}eG�� �/l�PD�� �Zf�bH�
�0�X��K-�9j���~�p�s<�ṌF� l?��51�x�J����]���//Jdܙ�c�@����S��k;;���>p9]�cE��K�R�o�p+(�rBr0��.&%9��5�k��|6'�1�=�zt������%����g��F�$�:����Ix+�����f���ذ���!�:�֌$�7®��Mh~O�#��3B�vC�%�\��1��z��ϗ$�}��I@�bw{���5������^ �L�rb���������l��&ʊ�TO��G�E�5\������j��>(�|����Q{0dk�V\���E�t柧=a�`���<�g��8!٦�G�˯�v"#�^�z�����e���Xޡ����	Re�kS�C��V9�w�g�ɛ�����+�N��%L�v}S���"3�`��q�R������x��0�U� Q��i�[MK��k�
�2�I[%%Чn�N� ��T��A?��ˋ���|ܚ �e��#�L�p�c�I_V�`y �:�-F�ӣL�^����^+����?���bF���4�
<��q(�L�t1��xTW�;G��<jY6z�6(k]�(=<xǪiUts���HX�`cè:*m�����2 �����b��M�/�0inǂ�2�5�z
A�_�x!g��ۙ�>ē5J� ��Q0�Z���e[��o;���M��t�E�TW�jmx�U�b�:Q����D�咉�7����}s��G�ix��+����Bc��@&@4�X�(~D�X1�U@}7�z�͏V��P������^f��ƶ��
�y�Zwy�[7�38U#�j�m�^���2\s��l)��H�u�Lt��}M��ͪ��K���΢���e�s.���!�O�hu6�5fb��kF�-v����`�!�S#W�o}��q�
�&�Ye9�ǔ�0�
?�MSV(����d��hc�ܠِ��Wŭ��b8U��W�d�t���3�+<9�x�ޯv	�e��r$ކ���w4r�p���"���Y�W˲�W8\�?\L1�T߶�`(w?@^��D}�^��lOid�`zxf-�5�kR�h�֖�ZHm[�jQ�_mqT�C"a>����,i2)#/;5J�V���z.�e�Os�=xf��}sl��'9������`֍��NrEl�B�YL�t3H��lm�`��5;W����q���ȗ�X�S�ׁWs�v��m�Iu��g��F�SC������jĖ=��{�;F�=8�_O�Q�\���wu�ϪC�cS���v���al�G�x�W.��[s�~��i��*�:�<w���n�(Sb����Q�>���9<�Y��	��l[��K��V�Z:��!+��t�|�K��|����25���R%�+��с�̋�9K��\0dw�/���8�	����n�ѱ�
,4E-�G�&��F��|?�j^]�w~'"��~>n������n��0#�fx�����t5=̝E��q&�^���TQ��cr��i�U����ח ^�E�,pΚAɊ&vVa�o�`cں��+���D=�x�n$�W�}7��=O�'Tc>e.�c^��>p!w�Y��v։�pӸk�e5����{�F�'(��5���2�Zi�O��g�t�-JsCs��ḼI"G�'�d��@�yZU����G̰������f�X���8��5�����(x*���y���mڴ�v�:�v��@u"B�.�؄]�ϲ\�9⢣M[Ǣ�v�}�v�ьZ��JhҖ��C�ƔX�7�K�i���i���x�}�HÅ����dP�ܑ;��B�m�,�0&zŵ�1@ДT��!*�H�S}x�HB��ʡ����7[<ƨ�F6�O,Q}���v���k���ʋ���u�j�>ے�u�<�
3�W���3b���aA�U]�A��ԝ��d�~,2�@�#��/�X��Ꚍ��p��u@,�*y�J�<�ճ���+=��PM ��_c>�6-��!��PW����6.���3e�uA�V $F-�	
_hx���̂ ]_�fq�˄}^�f���T�S�����ګ�H
Vc������A}̓\�3��*��SH���4��^�Ƭ��*gd\+췊}>63 ~ �y#5�$!�O(r�|�%2J|�1�u�u@����|4��B����Z����xK��S�rK�@l�c\,�pO����~�f��K�3�����S��� �Xէ�R�Q�Z.��s���#�⡭���5�T*:�A���}����^�F*�TÞ�,[(�C=��+"�$�9V)��"�Ū��Q���T�9&�L(�c���r��6�=��&2+��j[
_Pp��Nht7�;�WV�>;��>6ϰB��