XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:���ag(x-?�{���r�c��%c��2.�rA��N=A�@>�ߙ8��8S���zΔ��Y��-DR����^y`d�sd�cB&�m̊z��
��*�Ը�c5
|z��G��M^��).�2`�=o�|$���6����Hp�����/vM���۬YI�l�hK^:�\=�B�Kr!�rc�
�����[���#��~�'�U��J&y��ujp=k�$�F��l��O�1%�cq�����~��g�hM��U���U�.n���lH��iB�����6����y ?�)֯�s$�m�S��"�*��[�2 ���<CaL*��'m�B���ka�袏��7��y�,H2�=�̠��i�Hthnj�Y�;��+ʙ�(�XWA��mDI`O�*�|�p)NH�N*�IK�HA���ʵ�׌r����̼�kY'��Z��������ł�[�cϿFL���t~'�_��1z]`�>"�ƺj]�������3�GVʐ_Z4�=�����>���ZȎڮ�3�������u9W����;YA&�.�%w�-��g�ީ,�cF�D���f����lۻ-49b��w�=1��1QIѶA��2�L��M^w:��]�7T�7�[�p�%�r��"������t~�o��$t7N�Gm`s.U�ٹ������>,�x~/��s���� �-��\����@ط�v���ɀ%�L�����Ȑ�uC9)op���Z;��9�s[����g&�� *�XlxVHYEB    9732    14d0x��km��m�U(8���Ԡ%�B���˹o�-�_9Pe����l��%x84���q��}�F9|�|=FR�a\ �y�k7�b�B2}���̰]Do���v>$�����V���w/��x?��}]tǼ�.��cd�_V @��La�y�ݯ��ݝ�ݮ���v�o@�;������a�J�p��k�T?��7�pm�ބ}�)�]���i���D���R��Y�m�bm��%�A@
-��Q�х݌|�8 .����f���[���]�P��zY��;2�!!������ٚ(�is�P`v��z�j����8y�ZkytVU,�������#)YR�e�-�q:�25��`�����3w�Z����Z���8o qD�CP�'��}���<����E��p��R��B{�k�x!Q[� �}X����l�ߢ痺/f1���"�$Js�'�%�b�n<���R�熽��XS����5O��}���i����8�6���m�)���*�X���"'dCz��7�����P���ճQ `΃"�.%��PY�ۢ^�8麅�Z��]�?��K�m������qϸÿq���9&��dU���3�.�4�l5ԽEp(�`O��YUk�>\Jb�/ �)8p����>�`W����qm�M�+7}oP$�i$�7�n���ʌ�~������\(:���?*���[����KP��Rb����nK�M �]�F��w����R� ��
�gQ_���2�rI���O����v���b�Pͩ؞��"�$���[��A.�1��B{��P��.1��v�r��7a��"���[���x>��'���&���&�斈���"ϲ�$�d�ۀ'_˺���28�"y�e߮��[x���j 9;��F6�>��=!����l�B+L8h���]���N���( ���U:<�N�͖uH���Z�k��
A���!�zz�[XT��er+ �q�~�e ~y$X�C��B��Q�L�,j��P�%<٣��f�\x�.a�Ӈ��@�L��:8_��B��&�ctt����I
��dx���{��tR�򈎰��Ms_8m���*y:	h������	�  &�O"<�@4T��t���ru����aN+�� ^z6}���cl:�vP�������]E�0�熔����R7VkϘP�Q�y5���ʰ�B6���!\if��&���{V�"�k��E �R�`T*�G���tE�����i�k_��4ʿ��Xu�� �8�O���<�H~}���Ui܆W��9z���$fvӦV�J���~�%��l����}���_�+i�`?5d;x,��yw>t}켪�O ��~�,�ñ���M�J4n���j��	kF�+ ���A]���)�����O0�k�I�ݯ#��Z�y��X=UW0x�;2��f�ϡ��2��Ln���� ��W��zʒ؇���ǀ�v3\�*���!6�����ug-��.�%���3I/w��?��-����7��"��Զ��z��w�@0��E�D�F��!$��e��i��<�kv�(�W'���E�'|c1-�*w��'����n��;�؎b��F��)r��i���F$$w6�%{>�Ug�v�8ݽ*�6d������e��g踑d3v��}g䯶�0����\SyFD�ܤ�}]]���(�SmS[���7^u���K2�&�]��L���QC�V*ݥs�`M�۫1P�w��j��xΊ-�k*nxL�#]�R1������8����j.#�ksqW�^�U�(+i��S������n��u���RI�r�8:�0�Do�s���$Wxy$�M�����Ph�v�0Do,�υ�����7�짱��ZN��4�#�ư-7\�pQ__��#��S�mhj"�����R`]�ȬX|�-㸴|�$��eǫ3����Ns��=�z�h��o�m
�����w&�j��EZ���Q�y��(ցAcs��\@�G�̖��`�{u�<W&�NY6[+����긨�&�t�Sd{��"��L�j�l^%NpH���;�(�y"Fe������.�w�x�Xݰ=��N�$`+}��<4f����۞՞�{�=�M;��NMf�:�2�8\��H�R�h%��+��F��//�a^�B��Y_���_�ɡ��A~?s���d\8_,1�G=�P����'/�#Z0�/я����������|d�	��7c��q]�&A=R��#� �C��MO.sM�^�Nv�e{��1KF�G�?��'��q{�m������"�G�~t��j�a�W���$�U8� 4T���zp�D�@�5��dfC����5���FF�隝�U��Y����&�Ǖ����r[a�(ş9e��-H�c'�*��Cռ�޼b��������n��Ks&���ݘ�*U�A��M�!8����g��e����Pph��x�ҿ�4�WF��wU�&�~$cB#�XǨ��Tubv��%ϡ��*�&��yco�za��;8�z��oU���"���6Z�^^��|��&sݻѸ�a��,%^��v�j��8��s��^Y<xN�V,I\����s�A%`)c� �O�
=(��`�B;F�AZ�v�|���Ovٮ��fS���O�Pz]`.hﰾB��X��9�_;Ɇ9.T�H�j]D@�|�x�m�PT�kePK������W��rn���>�Z����"�� ���m	m�d�!����OޙCd��J +qHE�ժ��cP�Ī!�����"�c^�I���q���h�� ��Z0��21�^)��eϯ�r��ݽ�B��c)Z�Rp���	5H��[�`�Ҥ�`�]��x��erR6ь�����mo}o��ƗSf�yy��0��<�΂�ڠ�-��aX{y;P�H8|�۰��Ї�2���0�K����q���Gޢ*�uᗛ�8�m��>B���gC��nb6Cc��T���x�8�=�g���^Y�R����_�/�%q�n\NI7���dy=��&AE���qtؾ	�SJ��+�24P.L*LE "���M�r�*6�����I��Zˠ�Ҍ?�X����N�[d[���|�
WtcnD� ��/��ύT��hJ)��a�|F���g{��\�Y�S�)��������:Dv]�=?>1�d��+&�R�x��Y��_BQ�Ě�&=�B���5��Wt�?����G�\h��I>}�[�sև�q�'�%8ê��M����)���1�����i�W�bؖ��נ-��z���	Q������J�b;��T�"�,�Ɠ`�b�M��+k����|��~#�F:����>}1�q��P��7\?�ra��TBv�t�ADq�T�7q���b���x��d*�.c��Dє�ɳ� a��W���o��
�c��1���%�D�[�� ��4��3��zhm��ӵ�ϼ�r���g����W�,)r���n�d��ƶ�ӷ��a��,pث]�*OW�{k��' _�q�6��+L�u�L�
 ����_���+��M�i��]:|���f ���}���xޒ�����r���-NT�e��,�OA�DI@�p�T�Wd�h�_� ���NZ����u26��۾ўC�tUrg���Y�_ۄs���X��a�_p#�fEOĲP�[D`�t��n*f�� ��<T��檰[S�V�"aǵ�t������P�_��+�В�]�gz�d��?�[��:y�r�u�PXV����y�����p��O1MO���ə9���%/��tr�pb��F7��λ�k�zZ��]�#���̄�X#K$�G� p�uA7��P�E��r�#H��}�H��<�~�	���9
CT�{��p����$��_��N��_5�͑��z©D�`'ol]���������tjiv����T9k~2����C�����Nx'/�>U8�JG��n���N�uK�x(tL�������=w��>�lC!�xf���W��_7�9��ˁYސ��/�;��V8��o�5o�+�"#7��q/�k,��9-�Ŕ�bi����w�o9�UN8������'IE=Yd��F!a�Bh�3����x@!��ؒ��V�r��\��Nj^\�ѽ�h�>*��e%;��������/J`
i���A�y�8���{}�BH���[����KMY���kB��w�]��!r-��0M��CH_����c��l'0EFF�$���u*,2��E��Rt84���,���B� ���S�^9ƹ�C�c�Y�C|���7ƿ�4���z����h�BӇ����Y?J��R6'�Fԩ�wKB�x�'JcoYg}��F2N�u�h0���@"L�?f�eq��В!ց�ߏ�v��pܫ�����'������W���|�c��M�Va�=7Ʌ��ʇ.�5���B������">��r��"BAX2'w	
�E�%�%��rS�f)EF�H5���D
�:�Bɲ�
�C������t��a�����߭�aiw-{/3+��9{�wT����?�{���%��)����|kЇ�Tю8�Bl7k	o`W{�8�����R����L��� �Uп$�>ڍ?�[Ar�$�Z�Ă� B�j :5�]-�#�>ao�f,D{S�S���k����{yl�~w��j5�{��j�.����	�0ᖠ����l�� �=¯w�l`t��`U��:�D\���wUHLpP�PD�`gT��c��I%�@�ߑ%��:Yߒ����1%�ĳs��
r�hqE�
�G�.�����ӹ�^���w�8�HW8[���*�.�cHAUX�|5���&mR�:�����9h��.\&�<�=DT�\Ǩ�E�d���Q�i����]',`�;j�4�x?�x�4"� 7Rg9�y:�gۑg˨��:�I�i�կy��;�p|�iHǱ��K;�h����{���+��s�����Fơ� ���KK�&Zc98F���	�X���Ѡ����Sә�)��uM�w�Jã�J��jn�~i��KcK������E)q(D�i�p��^��pa���V���{*�	�CQ��8��pãV����|�l(�S�Ox5�)��R�ʍ՛"&)J��[$���@u"1<F���P�v���xТX��$k�/~T��g.N{���2Nי����+aک/F�+dK�e� ��d����;h������m�\LӁ�zv:f���0'ϮesC^b�!E`�ʣDB��x�a_2�Vf�������y�5������p