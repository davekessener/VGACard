XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����߇fmz�R9��q�$սD���E��z����T٬~I������Q�Ox{��������Cr�y��\x��Wy�SY}吪?˥Lf�G�3���s����.L���
����k�3�_Dᄕsɝ���W&�F�G�j����5BZ��r�h�<a\��*jqC�dFe'WT�LWØ��\��YWʤ8��Y��Tn*�w�����EE4{��|a�JRc�1�T�bN�g��5�{�?2{LX]�ʤj_Z�QO�G^����;���Q�²հ"��P��kP7b�d6��띓�ގ7�b���e��C%Fh��_R"��7F�
�E&Mf��{�v����>AP�}���j����o7B��e��;���|Ǔҍ.%�듚�k�,��Yr.���ɯ�$hp�V��q+ɹ$�a�P�������p���0�\��A�A�����z3��	�M��Ƣg@D���Q#�bf	(]#����[�a{�c���SB��u�j��/4��Hb��q�� 3�=�А�q����t=�EC'C �;H�K`6�st��\O�����7�<	ݔ����56ˏ�c�Ep:�U�ݽ	Qd��_ŵ�vm���.dYr��/�*$.԰�xl���L�)�� .p"RC@iP�[��M�����E���RCɿaG�Ж*�t�н���ӻ��;����5��Q��&7�?S-2
߅);��-��"C,�[C��|�0X����y\���jǷ�&0�zN?X9����G��}�7=XlxVHYEB    fa00    2d60�<y���r���D���U�Ta'�����H�"��8�G�Ifk���aiSC���VaڟQP�D��F����dz]$x���5`�rI��b%M��|FN���E��*�/�?���^����!8L,��s��\��}L�J
7��Mb0���>Ļ�_@8���g��;M2����(C&���Г��^8�nl�r+j�T�=�n�v�!gn�Zo���e�b��I5��о��x�yM�Uv-�v�0�/WcG\vX��6�8�_��#Y✾b#s����:�8M~�xɲ��js*TW��O�F�W���/!߭8s8�TA}?
b���[��<��d���;A��vz.׽�v��-hw����-E�=%pH5\f�^��UH�(�`�%��$�8���>j�NK(@����Ņ�w4c+D�v��gǔ��o-$����.�5���� 6�A�"뵤D�x:�������\Q��f_e�D��[�)�${b�'�f����yH�̈́e2{����$�=��x
Y��/ȧ+�avi4U�w��moO-)�̓sq��Jyb��䇵���Z�O8l�&X��0`4�q���`�����~�_��jյu��l�ˍ4�߉�G�JE?�^��8����ejp�ۣ��dĩ,z�;0�X���$N�=V�5����^�s���6\�j	`p G�j�6[� զ�4�d_*��z���$h�=D�$I�eV�x���%�Mx�G��s������#q�s}��E�����ml����� ���g�H�{�^�$	ff&��G'~�K�^o�=1����?'�$���VR���Q�I�7[��$�G��j�wdk��䯁�&��|op؟�نR�@N���ĳ�<�+�j��lmu�J��~� N�����Bh�����" ����J36l�ω�w�<s�7�U\���ֺ��_Չ��դĢPy
�j���G�����	װ���k߯�g�.~=�(�S�r>/Э�u�^��g��:�2ՍM�܈��QP<5x�vߜ�'��
����Y����vF�u7�5�說$5X��c���{UGQ`�B�vy5�:n1F���]����`/n�N� ��.����������Yۦ�GO�@�s��&�fB7y]B�k.g7�hZ~��Y�7���Ю��~y���P�@��9��t:�R~7?�W8>�Irư2�٤�f��R���t�J�(_w��V�ڇH�G�z�.[�Q aAٹ�ɥ�j�O��5e?G��lB�AF.p�Y��2�d�ў^9ϣ���FU1}Eg�ך]��gz��5>KE�E�)�fz8g{���W\xm�H
�4{޷E����p���>Z��һ=N��E���N�Sx�I�}�~��Ag���*� �u����6h(Y$����G-<������z#�f���n/���c�	K*c�'��E[h�S�q�@_����<�K����[��[��3�����)��<�����p��׶O	�=֊�#�������Id����~c��kn�� [<�jt���@���:�Kc��$�̈���8p���ct�����vF��Tk�b��0�P]^ݒ�S��y k���y�CߑOXe 5F�Ц	��������gn�o��z���#�-��+H��_�
Г<�Ͳa׋�������iU�U�dQ�	|�߾U���$�e���P�����)mZ�z�@��i+J{�u�IMz�D��W�a��q��:�/K�ɨ�_�I����wR9���gLiq��z�b�jؖ�ɫ4P#c
c��\V�/���Qa����� lF��q����+���5���e�e�������C��#J
m�?��zc�+m��J؅{Q�����wg��io!R��Y��vb�ޅ�ҋ��
3<�>�Ș�!��;=Ϻ:���.�V%���i���K	<.I��A
	�����U~0�?������� M"^��ؒ_�Pzߗ��F���\A��N�7�}�ep5�ɖB�=��y����X�~�$ �V�ƹ��v�D���[ �_K��$��=�����i�T&�AlD�iYxew"���8��$�.���j�B�A`9��r֡�W�j����|.�U�H}e�����3���G3���G��	�s�~�����l�4;��I�y�IC��5�_T�C����gӵ%ZI
�N��48鸀���!����6�j�$�0�����������d�P�5v}`��,��Lط��[��*V2Q��<"Xp��ʚ��J�y����qR-ŕ�#��<�4�!u��MS[�����7cȓeܩ3ę49�¾�*|���Pa��"Ax71���7B�Ϡ}��~���w*�hp�x��Z�ۘ�.�u�-%B+��#��~0�ҘS��� �i,ֻ�(�u*�E ����ˆ�["0��˱:
��<��/�Я���pVH��T��l� '9���al)�n��/��b���,�T���aŅ>X�JbP��]ִ��n�j�������s�[R3�u��`�@��@��M-��s^�B�C}Zd���y���q͘���Fǚ�4�q�+��F\�J�#���0x6�0����u[.�5�V�Z�A�_�e �V@~!�\ ��	������=qXQ ����A��/-$p���raZ��_��^�r������i�Ļ�q0" �\
SUtk�nYw�~�rt�U>"�9WL�#
=Hk��GU�T����ϟ)�R��Ѧ������ή`�[���9�Z�_�ޕ4*�U���B�M���J�4��mv��ZS����K3@T��xs��zGih�:V��1٣��u{��g�?8V\�ޘF�N�P�~jL�#� _6l�$b ���zo��b3E/�e'�Uh���텵��WK�`�kؙK��6���i.�.^�ʱ����� ��PB���DԩBLꓚ�q��H��ʟL9�E4���o8�-!�7g���XV�V�
�[.����t��p���i��Ŋ��ߥ4��u��!�0����s����
naQ�T�0������ؒwǄ�TVJuD�P�G=��a�E�C�[ݨ�>l��l�����Ck ���"n�$��q�7��}�PV�Pu�V���v���]IOϜ+�uჀ��d�v�0� �z�!-� �M� 8�;� ڳ'��F����q��TwK�)�X�n����M��[�m��t�=�Q�e³yLo'��d^u�>"��O�yh���pTDt� 3���~2tZx�"�.).x|��]���f�~��v�"}|?A�SJ`���u� ���*,S�ڌ��P(#�����S�p��½<�j Pt���\hE���ir�NY�Z�u^0$�ƨ�-z��e}�o��Ѣƃ{�Mi-L�9�׌��D�}�F�hl:� aX���*n�����R��IA e)����[�i�Q'��X�U���%fHS!���j �{�o/������g���?w��S�Q�ZĬ۠�Mx��W+�s�ׂT�W����KQ$4�������QUƶ�-_��.�ed��?͐�C=�;�:=I]-L������**8���P�'��JW�����5.i��2�V�o�f[o��(�+�K�hLJ�ն�W�~����f�i+E��7�vu=:�^
�k�^�1��}ۮ����;ɨkG��o%E�[�A9r��alȩ��t�0b_�Y��"<��"�@���*Uh4�)֡H~�zb�Y����롞x�*�v]�O�I1�!Ngk� �k�C��le���9D����밷-\�%m"n���q�Uk���̾09��zm~Ȉ�|�(�=��{���f{��]d�����	KPpVt��hƅ�Y�(v
�x���g�����>����sMo�$�ɐ�w�Q��@J�� >��+�����{KM���^��!v�dU��M�G�1a��3~�Ûa7o�#�4ԛO��<��GcF�K�/�!kg����r�ً��۾O= �,��0�SF���'e�7t���Wxzt	��a�:��˸��q�l�-/�[�� ���ln'Q�T���u�����iqR0���F���3�B��)[�i����V�,υ����(�N��i����?��wOh���)Ud5?��#�kB=���Ҿ��f�s룟��V�ze٦���鳉krXp���'�G� �<廨~2�̗��{n���?�����&0�1�m�E�'����_�(�UO��bk
`4�}0���u�P��$z��׆)�h\��q-���{�PF�q3N�`>�|6�k��B���;�A��ΤX��)�=vg4Ǜ����B��Mˁ(��WЏ�BK������|��<�R��ޘ�J�����lX0�x�n+�=�\�m�9_�Mb�0���3¼�-H�}Э#c;̽�T��!�Ib����Ԟ��fv��}C�5)(��1�}��%�xŨ�Y�Y����� r`.�X�����8HR�]=N�@�:��u��qUY��zJ��������: �O��آ��l�^�䳫��z2x�[8����@�����`��R�)�k,�n�oT�ך0�t�_�L��Kԋ=z룝����_"�Sù�B�-�2�H�l]�!FJp�Ӥ�r�����/��\�g�J���"* �L �kTeOq:�ȭ�T�L�6�d<��L�M?�'v�j��b�=)�:[U]]���׸�hJ��h��ngq�[��
$H�S���t ���_�9�	��xm�2b�����O|�Y��'X�>/�\�qU��y���\-/t�����(>Z!k�a7��ϼ�h��t�^�.�Ŝ�{�{�SS}�T�i�d�"~f��Z��Y&0�,My��;M��9��O�v(���QܱX���őQht޳�"v�J���-�M_p�>�kd��u�q��쥀6� %�
��bD��A��<f����N�fK��=h���/���Ajwk�l���Y�s��QK�H���Mr���~�<�����"�]�����PUd�`�=X�krF�
�ۏ$��Z!,�#j$�4�r���Ylz��>.T�ޢ
tN�J�ݽϯ��H�w�  _3Qb���%A�VP�QXS�L�c����n�V�lW�"ս�C�����+����������nΈ�à(;j!�ɩ�#V�������X�VS����.����X�a��|���|�/&��~U9��3z��)M����^(�.lc���7F��|��Fe{s����p�&�JV�Ξ\Or�gL+�׍]ז�@H�2I���~dW�p������V�t5hl��M`G�:,`���W�N�e��;;ɔU%�lW��a��*��E�q+�)b��D%���;�W��V�jG�h�b����˺B8fvD�é��iP�]9�SF��� �ɳ+��Ln�i����鞋�zwa �ՍC����|�8%���4)ǯ���?̐����}j/v���2^"�#�]�۾��z�Ίmr�s��^�C/<:v��U��T��i�6M�4<��6
#�)���A�Msǩ6]�n�f�� }���7�X�9�Hje������\���d��!`���	�`�|��MF$*��Z�yQ�ݞ�-elii9��$�CхA�cU�&�������l;�&�Sݎ(�N�$kR��8���M��mˢ ��ЅG
���k H@�F,bnI���|������ʩ�2\�
��QºB���<?��� �Fش��=�_�����[}ԟ٨�޵m_s�4;��L�IS��D��bii�|W���p��x,�z����DX6>�/q��AB�m䈏�K�Xyҭ�B��LU���+��
��6��~�i�%ӷhHghz�`���Q�p�>,�8m&�wZ��?�T�S�t��X��Uv{%��(�`&�/��s������A�W�(`�?�!Nh4����#��젦�Ձ�@���[	dp۪G�e�|���<xkϻ+#�����͊�{Z��8\7�f�TGéu�<~D��]:���h�Y��9)�N�:�H�{ѕ�"�c��w}�y�g�1B�zP��f0�q�[����#}�"��$�(��̸R��}��`��\�����T��J����{�ְ����	})�g��qW��V\���9X2�U/&��~#�RE��,ʿ�I����)���h�џ��R����y� ��- ��A�;������l�	�c�?܌�]N���H�Kߑ7:������E��{���Z�0ҕ����}���Fh�B�l�Xq�fѡ�L�F�{�d��U��jl a����|&9�g����Ň�)rUu+̓�r�5"�p�a2P�-ބpI���LR���2�����q+�Hr8%�N��uxN��0���j����ޮ��9s�;?��Ž�����A$Z��A�����ū�v����������%�X5��
��j�W��|d��ڲ�Y�Tmy!�>�iGǹ^G���ܔ0�{+BZ|�O���v�ﭐMأk�~<,�p����7Iv��G\L,�=q5������ɓux^��~F�.�ܓU#�!NZ��/��� �������i����i��9��WS��@��3��Mg�\W�
0{����ۘ1mt����g�<�FG�=�C�'M�lz;��v�(����!�=7;#ɴ�0jDܑ+i�HA�!O]C���R��O�u�$S(����`�x������FZ�{�"~�d���;8�^ȡ�z�Wm%c��V[o���?@p͗anR#vz�� N8A����$���+��-���%�� 6�V�I$0�ء� u�l���͠A�����<R�㙰fL�G��!��BKP��J�pt��b���^�n	�)�'MQXwa���`���v�A:��6!�Dl�#�SБ�mh�Y+�K`
�<!=������z�a��+L�1yծi�o�'�`	�QDJ�En��ޤ�u�hp�����!2�1�z\р�k#l������W��۹[oI��P�i����cYE�,�燖��KMy"yI˰���g�U�)��~VdjϚ+�} ��S���P���o'���<o%+��(�PGS���EnF���<�9�"�+|�G�H"�2��!Kj j[�@�(�^`�N�E�����֚��m��3ޫ��ܹ����K���6T�C[�7������Q�AnK�P��OA����j:B����WO��q�4;��w�қK���b��OU�^�5zx/��M^H��&iIdٙȧJ�QnD�n���şY7�-&X	�)�,
��4/�*5-p���p �/�J�v���@V��N�<M�uc�ԐA��,�g�*z�]j.3h�M�j;�L7�I�{��d%�O�Ho�5�
�w�HG�#p���6�����?���[��N�=�
L��_ƙ���O�
�G_���F�����~`|���3����x�l��,s!�x
*@�d�}���lQ�3N��<�f[Qe��Fd��{�"b���m�:�x�8���%T˓l���e����Ǹ�p�1+S���=�?�	U�lV�q�c���ƣ��*�Ε����m69P��&�rXwԀ�Y��)��%���E�\͏���$TW����	>qҵTڂ\����$��ʣ�룞9��'�DF7�S�.EmSF	Z�?vjEh�`�|������T;ܰ�^��7�\�3kn(|ݡ�~�`�:���ui��,�(�}q5�
 �f<�Q��?�4�������3$]�S����Fo��]�e��E
�گ\fm�ݍb'�5U���4'	ư����,R�`�Y�� ����-x^\���b����3�B
���ތY8;���,*�]�N��ӴCn۔��7.�w��g�z�B7n����]��f�I47˞e����ynz�~yl��ߺ��*��DW��9�)���x�P�鞄�����0�[D�7��)�z�S��j"hٴ�.8�'����Ž�*��C+[Xم⼕���!�B3������0�������2�>v���3y�xsUݶQx�ţ��\��T{J�B�xMT7�}��h����j��:��A��l�ΠT����i;�f���;$���SH��^�$t`p�9����}��E�f�Rrx������;�G7	�w%a�;~�{	?>��9V~�?�FS"0��򇂈�p_��kC�lT���}k������`���$z�����ՙT�kU�,mdZ�dǅY�n��h�ߤh��O;�@)S�JPL�T2�ɵ�-y�-����)�џIwO6�~`�[XS�v�sۓ�C�!\Ōot�ʖ�nWd��Uɮ�;f���Fo6{�7\�T���i�q#do��A�|���mmN�a<� �mp����m��=���M������Ri�]��=� |�͚�����)��X�=���,w{HE���E�jz�zˏ&_U���)ڔ�ʬ1F�+0<A�"D#�ߍƒ�e��v�,u�a�`8y"�;���Ȥ�������k�[��xt�;�uw��#f-6�9[{�%��z���	�Ѯ]��p���Ǎ:N�p5
G�Z�bo`�=��#�6&wB���=̻�����+M�7�yD'��ӛ/���gK��T��=\N>��5�p�iZ�c���������ɱQ�H~�F�NE?]�����!�m����B���*�Հ���t42�d}���]����Lu�X�7a5�S�w��8x��.��k-����P*	#NPv5�~h<�TȎ1�m����˕��7e.��ܘ�3��k���BdP�I��g�\���h��cHEY�������6B;���r2v������^��u�e�s�4�wp����"j��i��\O���r�W��z_gAՄ��湑��4b����8�%�z��U<>�g��&
��U�I�U,aC���"|1n�<�U���#�߿��N�Ic1��k�����!�&��9uE�pe$��V �a[��y���EK��k�^\���k��8�t�"X��H!���Q��?y��v�p��lr��Oj�ttY�v"Gӳdn� E��gP6/x5^�^:؅�s�Ο�tϜ:$zsU]�;�jhn��ѭ.1����x�'��%�#breQ�Gt���]��~�/�1Եk��Q�;�f�E�k�'�6�i=N�]O�4v~/�H?��mЙ�Zb��y�%1c�p�!��K�N�'ϤU������m?����1P���Z_�.�	�u �8�x^���yG���g,D0%r�f��?��KO��^^�Β.��)��Q:8D��B�'����Hgaf�ө�q~��;��8�2�u�*ޓW�G%���8RXՐuO$-��(t�$�7t< ����&�_.4d����2�#,���Av�OT�6�
A��p_$|)��B�W����Ô�0�j��,���O������ِ�>#ɜ��&�{p	ݐ+�c�^�)�p�ÂV��9�L���X�3���YEю��0�rm�S����n��ϻ9�e[i��~3aMe]��
�ɕ̱�������Q[;��)�ʡ��=�1Z\�M��-Ŀ�
�F��$qi/&$�ϟ�I�`y3�E��l�B��$���	]D��U��3�� t}��Q��󙶵��J�k�������-�膋u?�h<���sP�Kʠ��X��|e�� es�����(%�nT,�k�j$���&z2��h�-��P��~�	��S��4^�cK!ޛ�v]��-w��/���uu�c=���w�SBH�|�SG=��#�b�G"w^�a���mh�ʪ��� �����x��/d[�_L=�ޱ�w�)�o/��(G�C���j}(�����.���o���i�Wxv.@$�J��3��j<J�&7F��*��]�XV������^��|���jI�U f[�/�B'�~,���&ka:��5�7ä�Ԗ8��13j�y�8��Ch��qJѥ�/����O�P/e���9݇J⾇�����!c��;�=���x��d"eC�s�M^��������/��!���ƣ��|��� �Ѫ����hͪ�H@.nl��	!�0q��g$=�x�E���2K�6ǵ���T�L*�T�/���W٣ʫ���_����T�ם%��0����v��w��6բȞO�^<ڡ=�bvFt�{�+"���\�p�YH��I��O�[�������fK�#�D�o3@u-��\�F��A� � U���
ݩ���Hn���@>��J���J�T���x)� 鲿��3 ���|��J��s�i>���ii�D4/���7�c�8=�29��)�͕�����o����)�>���Q&l�^��&�QA}���`/4.U�3���R��7
K{ޚO$���_gp�QT`v��"��1=�Ǡ�[Z	:�0�1�b\�FǓ� tN|�9�̽r�R~������0F	��0�hy?�>R�>t!2��Ȏ*��4Q	_�5��=�I�(��~�mj=U�f�G����'���?%(0������ ���#,��Z���w?�ϕ?a�}���P�S�w�ξ�@_|^i�m���,�b1�x���
}���C=X���Qٟ��o5�����R���)Mצ@�wn�md=����z&�����KK��6�Qp��o���œ�s]"��W&E�捤�P��i����U"ϼ������v)g�i<��m��N�%U�� x(�3C�A��-T1��a��5`p	u?��p) �kM�E�{���Ef7
ۧx��).f���755�N�T<��1��_�+,B
��b���~�T5�J2's ���@���C�5�WB�������܈���VY-p�H��w��(J�y�X�j�H�(�zU2Ut���{%��J��b!���V�[�	E��ٱ���v�bl�-Ҙ����y����rs�{9�,��fr�#&��HM�����0]7#�_�RDx�:RAۿn&r�H�U�W�5���=�S� 
�z��BI�8�����}J���6e-�?�1A�d�N�X����g �S'_����֋�+i�$4������-�@����ǯ -0�ﾤ��_,2"%�"�k�Y���g8wުEx5�=�����d���#.:�P#�H�G��T��J���Z�z�9E:������Hb��pO�NpD噧�ĥd�շ�qM@�F9����%ѱ�BU�_4Bt.�R������% ?�R\A}��:�>
m���'�o
�EI(�5����\���v)�� v�i�d���_�4��Ӻ�ц&�Ћ�S����I��H�қ�'�q1���+i�#�[�Lq�|�ឮ�^�Gd���i]���C��w�l�d���fAE0�Sv-���R?*؃��C�'q�(�BH1��K��ʚ�ulƨ�'�km���-��-��"P����Ԡ��Y�o,�S;��YD.��(Rde;�T����~ux��:y��M0�����$�"�3O��C��B8XlxVHYEB    5914     f20>UV��0�.-�bh7[�ځ��!�qA����I�E�����v��%�8TR�9��ʋo���n�S�W�zR��m������1:�X5�r��(.��"�R倳�X��WF�*���!��t�p��3 _.(���Ly��UvJO���@h@����&Mٕ�%Oɰ���S �� ��s���fB��v�m�֩ן��G�؏�3�;�8�o�A�D{a;�M�w���&:�k���.ar����V��/�1Α����S�k~��kz�QZ[�FM}�kvO�Eog��j���#�L���[�J,̢/S��qQ�k)����M��M��V��/@�c���9ꤒ���=j�7Y�Z�;�J\Ljv�w�>ƜE⚘�{Z�(�)�2��p֌���kM��?hGd�]�轙v(Xt+�� ���؞sT��I�+�ټdz�x���.��y���Ma�@0&�Ȁ
8��i�v�> bFg�������i|�5��j�̭4�>����+Z��
�7 �ֿ͘��\OF��^{�3]<垈�����H�x��t��V�.��p`h�3�ޫ����++��Z!n�R��{{���5J��8/U��� ��̓U�ViPm �0�,c�1^d5�����?��:o�_p�'k
�J"L`��sp�)�4�� >���k4�Vχ���Վc�xn��\'�%}���
 �6�ܳ,˿<*̇��N�ĿDp,����z�7�Q�!3@���a��z}�L<�J���W�	N~�H�AŅt$]����e{.�1��Wj1�cm&%�����-#�}�,z��_{�ܐ����!��{��kiY�����d����*Æ����i�R��D�-�[Q1Ѝ��Úb*�g��#�a���	VǃvQ�R��Q'zƟ[����}�靎�ΕU�=E�\�� fܭ�Q5u6	�(\�5�d�D\�35���_�n#��I�~z>2C��r�
� �喼_.~���B�^#lRVb����� ���B|n^c�c�	QA��r-��LV�����*S2��+H���s���EY�R
熘�<2�Fj��$�ⷎ���Ȓ��־���I�5a�x�nI����7��WW��g�w�h -�g"<,o�wA��G�v����>�W^ϗv���@�I�+�~Hh:D�E���ƪD��,�9�AF��K�u�`����B�0���P+.�Pn3A��I�w�7�"�oh����De�.���u��D���C�{����l�������]��i�eg��af�׆̏#�O�ԖǮ�b�}{��C���l1ڶ��~�����"�{h�k�w�ͤ�췑���Uh(��u�M�����?��W:a�7���)�nn����爰���[�OU����� D{���G�Z6T�����<9F
]U�Њ7DncY�Z�iX���X���>IgQ>����#�r�l���s�#	d�&��7!�-C(ݿS&*��i&�%&�uH~�*�cW�;������R慀?��)�~����v:2[����nHz$=�>I9�T_ѳ]�����Ԡwth���ކ���Z�YPX,�ګ����-Y�F/���p��|FOo[L�f��hN-�v�F��1ӯ��ֿV�r!O��c"u�ڐ�\F�ε�1�*�P����b�W��N����ǃ�0ˢ��9x8�׭��\xv��|����n꯾V��mU���Fp�*��>EC������Y,��|=<ȟ%#Y���Qe8Nw���'��\�[�B{���t0�l��U�I:h��@�������,����sN�f�k�����������=f*��`�F!�X�CHn��$f��Qgd�*T���1��6	!���2�b�q�������e����{��:r��^�I�[�JN�l=%D�,��ς��;e�M�����|0���V��Ұ�끐b��CVjX;]o���2�����}���~���1����Պ�F@��NP�w�S�暓�c)�����3�S��C�~4 �V]a�l��`��:&�����I���P٧v(	��y��켆1�ѽ�mi�>,�ԍ@�����OVC��[W��\�� ~*X��|-���s�~4 \E;BK2�N��g��]E65���ρX]"_�#�!�.>6�@K��7�Px@? )�lqk�ֽ7�Մ�M�Y�?Tz>V	Mʷ�E�W_��i�r��j�k�B4@��'�'5J	s���~b1�?%:�.���,�O�$��>�25�������$L N=$!�E���Gǫ��c�i�XL�4_�
����	��n`C���Rr�1|x�dCm�|��B#0|Bd�Ӡ>w�0	uK~j�}z���ɷx��� h,G�=�Xm���A�ʚ����n�8�r�%|Ǉ�?���x��@���ߘ��<����(��!�]��)~z���X	�R��O��te//"U)wF(��*EEE����J|f5��iج�����R�:Qp5K) � �H��I�A,l[q�~v&e��tu�e|M�(��W͚xф��x�a��\�X�P'��>/�����̓�{�i��5���"�0_� �eлf�CA�$����e���짠��,F��ͳ��(��l��C�T�{(׃b.���N�{�H��Q�U�tZ`M�ܩ���� �|��D�x���-|vB^��AF�YH����s��Y��y�|h��0�Z�����i�A�p�Y�K5~�u����u~T�xO-�Q��v�
zpY��J\|\/��<B��]6#�ޜI�x����8H�	S�(y�� �M%01�E�<����G��z����疵��th��L�;k����X�s`�ō��Z���,X��[:���d��C���O*-�#b��C�q* #���Vu���ZHm��%^о
�;��'{Ltjn{�:�J��>���Cla�E�3�C�{�J�E�'�=Mdp*����hZ<R�q�j�N�t�UFR��m�y(��y���hh�C�wh�M���H:����yNB���i�+z���'��j��{*���@x���E��t7XA��T"��5_WgUs���Y�d�zk�e19ټ��;3��Y.��UKv�p�4�p`e�U�u���R'��֤�3 3���d|��ZO���`z2�,F�6 #�x���Q�C2����'\/6	�	Rk�/�6钐����P>-��c���J��G�D,Ee�
��1SV3���Z��3�4��>r�"G�����ST"~�[�w��$��|�4�-+:Cd#z�D �֕;�����~A�@ԓfqG���M�}��k3A���;w��g�{� 8���1�"��Ւ
a��L[4�"���T8i^�9�N��9����g
&'8���Y_���6�U�ch�.��`�c���Tl�sv=��} �^w�֓f�bΉ�.���M��{�=����q3�ظ.�^�MUj����� g����/�K�F��5�zM�ƞ3���� F��������OY_�R��'��1�-#T�	&gn䥾�쁉c�ߡ���:)$�(���Ye���J�o6	F.]ڃ�j���(��]�h=��]�1�B�x�I��X�?ȕ-�OT� A���K@��O�s�����gbH[SHa�/��`榤���1�
It����F6V��++j8~�_q<�do����d+݌�i�=��\-��a[�6f�&�GI�]E%�~O����*j(�ν��? �����8<*)Ay�4�a�r�"���5�،��P���d� K�F��P��a'�
=O7M�0h�/��O��!�}��ٷg2Ѳ~�����c�vi-�ڌL�Jd�&�