library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-------------------------------------------------------------------------------

entity charset_mod is
	port
	(
		char_sel	: in std_logic_vector(6 downto 0);
		invert		: in std_logic;
		
		px_x		: in std_logic_vector(2 downto 0);
		px_y		: in std_logic_vector(2 downto 0);
		
		pixel		: out std_logic
	);
end entity charset_mod;

-------------------------------------------------------------------------------

architecture Behavioral of charset_mod is

type charset_t is array (0 to 127) of std_logic_vector (63 downto 0);

constant CHARSET : charset_t := (
"00000000" &
"01100000" &
"00110000" &
"00011010" &
"00001110" &
"00001110" &
"00011110" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00000000" &
"00011000" &
"00000000",

"00000000" &
"00110110" &
"00110110" &
"00110110" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00100100" &
"01111110" &
"00100100" &
"00100100" &
"01111110" &
"00100100" &
"00000000",

"00000000" &
"00011000" &
"00111110" &
"01100000" &
"00111100" &
"00000110" &
"01111100" &
"00011000",

"00000000" &
"01100110" &
"01101100" &
"00011000" &
"00110000" &
"01100110" &
"01000110" &
"00000000",

"00000000" &
"00011100" &
"00110110" &
"00011100" &
"00111000" &
"01101111" &
"01100110" &
"00111011",

"00000000" &
"00011000" &
"00011000" &
"00011000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00011100" &
"00111000" &
"00110000" &
"00110000" &
"00111000" &
"00011100" &
"00000000",

"00000000" &
"00111000" &
"00011100" &
"00001100" &
"00001100" &
"00011100" &
"00111000" &
"00000000",

"00000000" &
"00000000" &
"00110110" &
"00011100" &
"01111111" &
"00011100" &
"00110110" &
"00000000",

"00000000" &
"00000000" &
"00001000" &
"00001000" &
"00111110" &
"00001000" &
"00001000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00110000" &
"00110000" &
"01100000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00111110" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00110000" &
"00110000" &
"00000000",

"00000000" &
"00000110" &
"00001100" &
"00011000" &
"00110000" &
"01100000" &
"01000000" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"01101110" &
"01110110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"00011000" &
"00111000" &
"00011000" &
"00011000" &
"00011000" &
"00111100" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"00001100" &
"00011000" &
"00110000" &
"01111110" &
"00000000",

"00000000" &
"01111110" &
"00001100" &
"00011000" &
"00001100" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"00001100" &
"00011100" &
"00111100" &
"01101100" &
"01111110" &
"00001100" &
"00000000",

"00000000" &
"01111110" &
"01100000" &
"01111100" &
"00000110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"00111100" &
"01100000" &
"01111100" &
"01100110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"01111110" &
"00000110" &
"00001100" &
"00011000" &
"00110000" &
"00110000" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"00111100" &
"01100110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"00111110" &
"00000110" &
"00001100" &
"00111000" &
"00000000",

"00000000" &
"00000000" &
"00110000" &
"00110000" &
"00000000" &
"00110000" &
"00110000" &
"00000000",

"00000000" &
"00000000" &
"00110000" &
"00110000" &
"00000000" &
"00110000" &
"00110000" &
"01100000",

"00000000" &
"00000110" &
"00001100" &
"00011000" &
"00110000" &
"00011000" &
"00001100" &
"00000110",

"00000000" &
"00000000" &
"01111110" &
"00000000" &
"00000000" &
"01111110" &
"00000000" &
"00000000",

"00000000" &
"01100000" &
"00110000" &
"00011000" &
"00001100" &
"00011000" &
"00110000" &
"01100000",

"00000000" &
"00111100" &
"01100110" &
"00001100" &
"00011000" &
"00000000" &
"00011000" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"01101110" &
"01101110" &
"01100000" &
"00111110" &
"00000000",

"00000000" &
"00011000" &
"00111100" &
"01100110" &
"01100110" &
"01111110" &
"01100110" &
"00000000",

"00000000" &
"01111100" &
"01100110" &
"01111100" &
"01100110" &
"01100110" &
"01111100" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"01100000" &
"01100000" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"01111000" &
"01101100" &
"01100110" &
"01100110" &
"01101100" &
"01111000" &
"00000000",

"00000000" &
"01111110" &
"01100000" &
"01111100" &
"01100000" &
"01100000" &
"01111110" &
"00000000",

"00000000" &
"01111110" &
"01100000" &
"01111100" &
"01100000" &
"01100000" &
"01100000" &
"00000000",

"00000000" &
"00111110" &
"01100000" &
"01100000" &
"01101110" &
"01100110" &
"00111110" &
"00000000",

"00000000" &
"01100110" &
"01100110" &
"01111110" &
"01100110" &
"01100110" &
"01100110" &
"00000000",

"00000000" &
"01111110" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"01111110" &
"00000000",

"00000000" &
"00001110" &
"00000110" &
"00000110" &
"00000110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"01100110" &
"01101100" &
"01111000" &
"01111000" &
"01101100" &
"01100110" &
"00000000",

"00000000" &
"01100000" &
"01100000" &
"01100000" &
"01100000" &
"01100000" &
"01111110" &
"00000000",

"00000000" &
"01100011" &
"01110111" &
"01111111" &
"01101011" &
"01100011" &
"01100011" &
"00000000",

"00000000" &
"01100110" &
"01110110" &
"01111110" &
"01101110" &
"01100110" &
"01100110" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"01111100" &
"01100110" &
"01100110" &
"01111100" &
"01100000" &
"01100000" &
"00000000",

"00000000" &
"00111100" &
"01100110" &
"01100110" &
"01100110" &
"01101100" &
"00110110" &
"00000000",

"00000000" &
"01111100" &
"01100110" &
"01100110" &
"01111100" &
"01101100" &
"01100110" &
"00000000",

"00000000" &
"00111110" &
"01100000" &
"00111100" &
"00000110" &
"00000110" &
"01111100" &
"00000000",

"00000000" &
"01111110" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00000000",

"00000000" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"01111110" &
"00000000",

"00000000" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"00111100" &
"00011000" &
"00000000",

"00000000" &
"01100011" &
"01100011" &
"01101011" &
"01111111" &
"01110111" &
"01100011" &
"00000000",

"00000000" &
"01100110" &
"01100110" &
"00111100" &
"00111100" &
"01100110" &
"01100110" &
"00000000",

"00000000" &
"01100110" &
"01100110" &
"00111100" &
"00011000" &
"00011000" &
"00011000" &
"00000000",

"00000000" &
"01111110" &
"00001100" &
"00011000" &
"00110000" &
"01100000" &
"01111110" &
"00000000",

"00000000" &
"00111100" &
"00110000" &
"00110000" &
"00110000" &
"00110000" &
"00111100" &
"00000000",

"00000000" &
"01000000" &
"01100000" &
"00110000" &
"00011000" &
"00001100" &
"00000110" &
"00000000",

"00000000" &
"00111100" &
"00001100" &
"00001100" &
"00001100" &
"00001100" &
"00111100" &
"00000000",

"00000000" &
"00001000" &
"00011100" &
"00110110" &
"00100010" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"01111111" &
"00000000",

"00000000" &
"00100000" &
"00010000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"00000000" &
"00111100" &
"00000110" &
"00111110" &
"01100110" &
"00111110" &
"00000000",

"00000000" &
"01100000" &
"01100000" &
"01111100" &
"01100110" &
"01100110" &
"01111100" &
"00000000",

"00000000" &
"00000000" &
"00111100" &
"01100000" &
"01100000" &
"01100000" &
"00111100" &
"00000000",

"00000000" &
"00000110" &
"00000110" &
"00111110" &
"01100110" &
"01100110" &
"00111110" &
"00000000",

"00000000" &
"00000000" &
"00111100" &
"01100110" &
"01111110" &
"01100000" &
"00111100" &
"00000000",

"00000000" &
"00001110" &
"00011000" &
"00111110" &
"00011000" &
"00011000" &
"00011000" &
"00000000",

"00000000" &
"00000000" &
"00111110" &
"01100110" &
"01100110" &
"00111110" &
"00000110" &
"01111100",

"00000000" &
"01100000" &
"01100000" &
"01111100" &
"01100110" &
"01100110" &
"01100110" &
"00000000",

"00000000" &
"00011000" &
"00000000" &
"00111000" &
"00011000" &
"00011000" &
"00111100" &
"00000000",

"00000000" &
"00001100" &
"00000000" &
"00001100" &
"00001100" &
"00001100" &
"00001100" &
"01111000",

"00000000" &
"01100000" &
"01100000" &
"01101100" &
"01111000" &
"01101100" &
"01100110" &
"00000000",

"00000000" &
"00111000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00111100" &
"00000000",

"00000000" &
"00000000" &
"01100110" &
"01111111" &
"01111111" &
"01101011" &
"01100011" &
"00000000",

"00000000" &
"00000000" &
"01111100" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"00000000",

"00000000" &
"00000000" &
"00111100" &
"01100110" &
"01100110" &
"01100110" &
"00111100" &
"00000000",

"00000000" &
"00000000" &
"01111100" &
"01100110" &
"01100110" &
"01111100" &
"01100000" &
"01100000",

"00000000" &
"00000000" &
"00111110" &
"01100110" &
"01100110" &
"00111110" &
"00000110" &
"00000110",

"00000000" &
"00000000" &
"01111100" &
"01100110" &
"01100000" &
"01100000" &
"01100000" &
"00000000",

"00000000" &
"00000000" &
"00111110" &
"01100000" &
"00111100" &
"00000110" &
"01111100" &
"00000000",

"00000000" &
"00011000" &
"01111110" &
"00011000" &
"00011000" &
"00011000" &
"00001110" &
"00000000",

"00000000" &
"00000000" &
"01100110" &
"01100110" &
"01100110" &
"01100110" &
"00111110" &
"00000000",

"00000000" &
"00000000" &
"01100110" &
"01100110" &
"01100110" &
"00111100" &
"00011000" &
"00000000",

"00000000" &
"00000000" &
"01100011" &
"01101011" &
"01111111" &
"00111110" &
"00110110" &
"00000000",

"00000000" &
"00000000" &
"01100110" &
"00111100" &
"00011000" &
"00111100" &
"01100110" &
"00000000",

"00000000" &
"00000000" &
"01100110" &
"01100110" &
"01100110" &
"00111110" &
"00001100" &
"01111000",

"00000000" &
"00000000" &
"01111110" &
"00001100" &
"00011000" &
"00110000" &
"01111110" &
"00000000",

"00000000" &
"00001100" &
"00001000" &
"00011000" &
"00110000" &
"00011000" &
"00001000" &
"00001100",

"00000000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00011000" &
"00011000",

"00000000" &
"00110000" &
"00010000" &
"00011000" &
"00001100" &
"00011000" &
"00010000" &
"00110000",

"00000000" &
"00010100" &
"00101000" &
"00000000" &
"00000000" &
"00000000" &
"00000000" &
"00000000",

"00000000" &
"01111110" &
"01000010" &
"01000010" &
"01000010" &
"01000010" &
"01111110" &
"00000000"
);

begin -------------------------------------------------------------------------

pixel <= CHARSET(to_integer(unsigned(char_sel)))(to_integer(unsigned(not (px_y & px_x)))) xor invert;

end Behavioral;
