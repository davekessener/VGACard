XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t"G�W�]d)���6l���m�?Y\R�I���2t7v���
eN`�te9���4����D2ߋ	�9����hM��{�~��@H��gT��ȟ�&:1D���<�O[�:��Ւ����X��I�?x�h=��Zx�oP��#w*y��j#0�b����q����
S�*�k3-ó?�o���@�5�m3��u.� pv~}�@�ĆV�|�v�SnI].�J~���k�B���Z��|�0�a�rM��ºG0ϐ�&�M��'��,��� �CHu@�%�"5!�F�)�uw"�Jfy����/+��3s�b�ȕ��Z�(��9��*�Oy�<@a���"�:�3� `4?��!>�w�S��>��� ��Uχ���ތB��}ޗh8T�;��C!��!���kK��I�m�>h����8�ް�l�����5����G�|֍ۨ�0{�r�J��=���)
l`�H�]��,t�xh~h� �Ѷ��r��eC�%��H�i�W%N��)\}F�~�X:���M?
R�b�5��C��@��D�se�U�V�ͺ����2�I��� �I�۶{�Mq�`�d�S�8��sl�Tq�������p�	���o�w	��X�Ҋ��8M���:�(��X�ǚ���bt���C�~��݂�V���ʍ����{v�q�7���Г�5��\�U��Y[���N��C����vL:��hA�q���p���}�cR�j���i�=�C��R��V�� ��(��O���3XlxVHYEB    3042     c80���֛L]�R1!/^G�b�"��dtW_��9ˑ@�����B�D2vB=�A2b�8�9������z���� y�^ 2�(y����3�f]�]�l���x`k�qs�b�ё��W���7:�i.��؎�Ф_=�fOx��+�2?�㧭|
;B'�N��(Z�������V[��:|�j��y�cKR+���mBp�������2vH_�����ş�]���H���f���(�$� �Z3��z���Hb�����Etk�7����%#'*	�mH�Ɨ�z?�Z;:�E�#�g�|�t\�[Xb\F�
�G�����.��B$��kⲢ�6-d�vB��������h/�ct��e�3ч�b�%gaO���E�H��3��X�K��~���I#}j�sh��,���-Ugl+�9z��6݃'��V/������MF��H���y�8wŽ�^Fx��L��gg�3U�%3�
���be�x��t!�a.�o�K'Jv6sHJ�����ߺ&)C�
�`�/h9(�K��B�gRGg��$:;X�=�3�:)u[��eW���}�JY<�u��qX�#���]e���Yΐܒ%�M37��뀆5̓:��鄶$?8�C ��Z�G�pr��aClb\����y�A�%��i��?ª���*!�J\��z�RQ+E��ӪC�7�N˾cZ�,��},%����M&g��K�Z���/φǽV�%#]<���~��1E�c� V��e����\���<,{5̵d�P��tih4�iu��|Y]�w��5 �j�D��bg��@�o�������WD��跋˾��vA֏wcl7�S"#(���ա���(�8ge_*>Q\��G���d��?_���P�8��ę�3:�U
Ou�5�o��<��X���'���/2`���ûX����W�.9�vD�"��)��OU�Ă��j��O?�)^����?Y.iM�e*��(�dÔ�~�9骐5�^�y�R����g��&g�9.SVo.�<���'�.�±�������@K���V���z<>=0�rۼ�A^�����B�����آ�ü����,����#N 03�~��y��B�Аy�a	��'�<:�w��gJ��vX�����2��8�D8,\�������'B����>�?��`�A���ۘ9���U���%᱙��zz�/���l5T�e�5��ǰ}����_�Ȳ\ˠG]���t�+ȗ�1�8wO������RI\�	w��0��4�&���J��ABOa���p��B�����N��Sw�1o���G7��@0PN���5�v��{� ���8a��ߵs�O�(��Bz�=��3���X.����*��
�e=��66�SK-�7b]��Z]�=�$���sY�����_:�X>���U��
u"�70g�7�h��8��C��>�Kn���W������V\9_�'j���<�Os>2y���tQGR�ie��>�Y��yI׀��<r,ZA7��i�%�&dT��-	0��h�ss�\���罤K�����n-_�^�4��I�u����r��'����	���'��-	��b��Źl>rg�|P�m�b��,�Y���0%;Gl4)}���YB>�9vN��
"k翙���:��})��>��~*��{S���-� ֻ*�
,�j��\��9��J����|���ν#�5��X`u���<w�$��$T��!.J0�A���`�|[NԸ��#�<gB� �9�a��Bly�/��_���ZBR橳4H�T�잣-Z3c��[�nmV|aE�+��Y^z�Mc>\���& ~�j��'Rx��p�i��DW�~��40������F��˗���a�!	_����h�U����(�^��>��d�`�=u �2s�E��d'+n]¡�6'5�)�và^�Y���=�����m׶'%��.kk1V��U�P>��{�`?�`����:@@ɜH����ȴ���G��^��N�B��� =W��Җ+>=N .�2�x��-@ŵ<��L���B(�x���*����� ߤ6��4렝�>)�L��1�Q�mPX9?ϕ�`�d��jr9�N�_�Lc��1F	�*H\�)7��FʂQ ����I2�/�4lo�t�}C��%���B�_�=
>�2#d�C��O���iSI9�s1�{~ɁA�י%v7Tł>�A�kK�!F{̗xiGQ�����ω��r�̶ӝ~���Oǘ���3�y�6�;��l��(�+ل���D�.���Z�z�����]���I��5��u�}�ϐ:9�hu�S��֮#͡�� s/�a5ϭ^�d����w{��;�E��(�b#�p��Uܤ9��#?[/�7�Mq�[�0�❜�>$;�}[�Џy:�(�a�P|;�̩7����V���r���n�,	f�;9�����%��aK/^���b��>K�d0�[��ߣs�l����/�����q�����|���4pI�o�6i��rd.|Z��Zq��N+e>Q� U�^(��MU���Ѭ���#�}{�'Άa 0��q���w�d�N�p��U V��J�n��j��T�ﯬ�I��p��1�J*	S�W���RE���g�qI2en-�@��~�VS9z��s��ljDD6�;F8L�a$�``^`r�c!m����ٶ?Q��v3M�Va�p~/���1���֙�~_d Rtgm0���T�ǮҔv7^�5������^ >�+�-�KS�L"��_�̎��X����#*K�#2�)�#|�!��(}mV�.~!ڂ�8[��Z�M=���D�:ܵӀ���mZ(8��OI���٦Q�uA��+�����#ʎ��~�CD!�	�^��!Vzq4ssRٸt%;�7���g���1����1�b*)��}UL#5#?��h���ϹF�P8�OH�9y������b>�Kx~��oD|D}_�t���I�5��F'��[1U�aG�"*�`�^���t-yM.�=���r��qȎ����i����ڢ^��N��<o�M����|B�'�Iߚk��<��Xd�)�BCs�,ڦB����)fb�3v����XRҴ�7�Ф¾�0�76XCx�XgB�i:�D�����P֩���g�z����{H����d�u|Äk�=��