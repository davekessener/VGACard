XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ǘu��&�����׺�gx��Z�Tn<�m����rC�R�U�~��E3�,C����5,on �2�^xe��Bs���k̩�ɥ��QR��J[�I^�ehqc�#��	w7��i�>9� d�"8J�4��B�cJ?j�(݁���w���=b��S��)iB�K�U�J��L8�� Ej!S!Ke��	��`oM�b��3�C���I���
�C�(u�:��yѬ��SA��=T�W�cn�&����1y2�F$�'6���!kYf_|�[m��c˭�ˬ'��E�E�⮢�yA�,��d�9���Sv��M*"�^���z��waR G���{���ĵ�;f#���E޾��%67<a���W��6����E`�`�:�R���`�K��Ip�ɸb���&U��ۤ�QlU��G,��h���[C�Y�g���|��A��U@`;ͦ�w�7Sa"Dw��7�0��dQ�* �LP�F{j�d`Ա�����he>��ʕj�l�6�^rd�x)���N�Ӏ@x\x�5�.��H�K����d�XМX�bj�_�e��T���ه�P���A  �+.�H��K����D.{o���v'(�h�.ʻk���&1����;�t�i0_G���-�	8�o��x���,���{rA!�����p<)x�B�����������g��r޺g���c���;�� �SS���m�j��w��kl�DH�z�Dک���%EtG�~]��2�G8����|��{H6��XlxVHYEB    fa00    2950
|(64�f��"��_qE�'�<82쮽��+kW��]�):��e͍ݳ����+˕艫��l��BZ^O(VB��m}q�ڎ�2��i{o3�ĈXGETǍ2��,ک"�)q]4�&�u&�A	��>ԗXk/".�H���UUܞ��2?9�
������w2���X�&�A�	���H�T� C�|T�|!i���\u��76�8PC��J�O2��/����c�6SN1�����'�Y|�vZ��g�vj�Am������-����E%i��Q��D�� ���p8�?�`2yN�8Em¡a��y��4� -/Y6�b="��Wa�.��3ԯ�b7�1��ٺ�x�G�"��p��P/���I.(OW��E��YЄ�����
gɁP�-��b�@��Ŋ̈�g�#�1�xf�43Y��:�S�!RrpyWߌ<���r�HJF�Gӏ�E�wތ\is�1$]�:N���$-�3�>��9l��mJ�
���ko��Q ���h#�|��8U�,�Cٸ����T��"�)���b12�V�֤N��Q�f.���ltk�ALP�΅ ��:�lt��b�j�J_�+WcVB�4`�-T�0e�hQ{�|��`�K""��YhfQ�W� ���r��Gr�̋�=D3[j���)d�^���=$@,��)U����7:��Q��C�3z���$ϋ	�w�9�q����+�`��0�1o�+`fvv5|���R^���5p���������H�0���>�gj�ckb�}�+ D�Qm��}�͈�-��E/\~Zэ�Psw�3��_.2Aҏ��f�\m��7K�1����U0��L1]S�F-P �P�%��Q:܉�8}���as��@��Ʀ4+�@1B=��=�W)e�X�o&�����wWZ$8ۄ�R�#&~V���iwQ���xܻ�Y6Z��د�Sm���𖥡�	+��R�(d8s6й���)Ԭ��/�D��ukm�x��w��%k`(<6u�l���48%/�r�xq��\COr?���HO��)�1�]Qe*e���3P��h�O���9�9���tv=�+�0�˻���������,����}x�z����6���4�E(8�d,��+�PZ��WCZ�q��ǅ(=Ni<R���[Y�s��� &�өƲ�Ƣa�z}]cI�l{oAx��� �?IxR�g6�VV/���xɾ'��Vn�w|��]�0�X��{IK̶�^�^�c������6)�?'��Р�&}�<��6}e�+`p�ȫ�p��:�����`J������yƜUW�P��"��~�m��N��8��)Q��UݣA>HX������)�%�L��=�;أ��z �rd�������",$1R�+ͬэ�{_���ZH8�凐��Էa��Kx���1���#��<oaevB���
�:� �G>��.:���c���Z��W��aE����ҰK}����� :��U���ꩄT}z1��@������ຝ�m�\�(����,�m: iĚT'�F2B����|
�=4i�P,�&����T�7P��pi��ѳ��hZ]�9�L��X Tp��T��E7����!�q�h�'~�B���e/14���c$<b�s�\��A���{��Y�t���s{�y�
6��<��Ɇ���l��.N�afR��j,�q#	������oX��.�u���G8�����$�_Q�k��)��_�V� �g����P՗�զw�a\�Xr��n'�A�{�Dl��9nG{�7���r��4D�,���-���\-�k�CH<�s������up�^͸αn��V# H7�4��@H�uOp%<�	5f���%��LL��G�O�A�Q;��F=�)��_z]��#���ت�$�����Kk���_�~�E-��.�sl����?�Lv	6?=�����R:�&������XZ� �d��*�z��ط�Bt���c`�L2��^�r��>A�g>}XJ���X�C�?,�=�
�"�}GC�#��D "�SnJF��i9z�Ar�`��Q���6���.l�B�1m��a^�ɓ��)n\hz�)#��ǡJIY�u�9��,	��V}G#��G=FZ���/���r��E��8VҮ�(���0<��%#2�A �w��R��.-O۲[�渫�>��]dH@.��,케m����oX߶ZS����w_��'�a]\���M�uؗ���e���W$!W��P��ˤxcg����w`�|w�}|L�MOD���m�p_u�lظ���E�Dp̧��T��ZA6@��**!y?A h���J9�$w����p�&��"ͩ.[�:��h� ks��v�P~\V��L��#��تLO�N�[�QQqEgy�"����0�V��K��<q�)�=�r=�>�7=b�� RTf� �Ynn���a��0�MM(3�~��<C�Yp`�J3�[pJ,p��S��AS�Bj<�!�Q<�woAȧ�� N!�ܚ���I��J������[���	�ɛ���?��#c�o��8�	4�&����n��\p]f���s9��<iㅃ�p��I-�U�r>-����v�Rjy�"LY�5U�,¹x�.�B�!I?F���2��P�sk��s��R����$�6�J�:i3\�xi=�U--���L{�zz{�X�?�Q��k���>�ͧ+����-�i���+��L������xј�K������������T�cHSw����E�=�$d`�&��#
�˾-����T�{������%X��rnZ�X 	������_����JAGۦ"�-
䃸8�o�ڹ��6Pr�W#���� 2Kw9�l�����{���FWU��s%,�Ѹ��¬��>�¢6�/���1aa �n^p�+C���3#�����fux�>�/	D�������.ZݑHr�ʁ*(J������7�v�V����P+l�v����Dl�th�2���I���� �?����%ђ)�~Fk'���ɞF�̱����,X`� �TE
�V�7W���0� ���_ڍ��^�����<�yP��?X	�g �dʗי=�~���t\t�:�sP�߅��Ԙ]��g8�ݔ FVc%��_��-�}�/Pc��w�em��/�W=Pw��Q��W�SK����R�4���oS�#���VR8!�Ky�jE��x�Xo�<�P��cw��~3Kِ��l���=���:��3OL�����z�M>(��'�o�CN�LH�ְ�1�uN`��� S	BgX���'\���Ĥ��w�zC)��D�pŢ���)*����pM�D��xb6��U����B�g�8g� ��˥���\��x�Ϙ�k{�n�P߭`��Y2��ሂ3��
�{����*�T�1��ϛ�8ü��"���K(z��_��t�e�w|(�iP��e�'���!U�D|\>���m�c�
4�g1�2�򺫖�;��X���rR�Z�Eu�?UĈ����\[]��h�	%R�դ��EEO�ƪ��Я�����\��h���`���?d��ͬM@��B��!������	u���Acm�h�Db0��Ѩl�{"�%�L�.�K��X�1��	�c�?Bȭ���'���b�=�
�Ώmi��lD����v����5ܣ��k�\��V�����p�_����>���;2[�6���nl�ڥnV�ь�9�Sb@�>gF�]���sՖ�������ӵ�+ޚ,�@�FF|_���I9glhv9bG6QhF|��P�vK�u.V�T�4�O/��D"��gi<�؀�B*���ŭ�U���8�4��ˎ��B����Lu��/i!B�����;��D������t��w2�N���e�漜>��_ec,�CLe�=s�D�Ǫ��K@���"�R>=�uO�bF��#���3�^G}��<��d ,��N���ٳ{R�h������F����iԊBI��}mr%�FjW{Kp�V��h�\Qv�}g��U�2�۪)u�7z�2x)Sx<{��� ��y
~���4mWa�A�[�J+93�����}��l���d�%k3_R�~j�>�Ô�>^6j����{5�N@��U%{q4M�*� ���i�"�n�yY��yO6��
�	2�F��J����3����d'^yIX)�\�:k쒛#m_~\ө���k�t�����!V7�f`�pg�PIOv�;�n�a�����(_9�{���4$�hVZ�����=Ł���>K��,� �+�����">{!���5���7�h��L4�39�����9�	�];�R��h�dV�2�ct8'{8�������[�V�n+��z���5ř�!���]h�h9T�ʔB ���7.�ϑ�9:c� `'��z[��teJ菱N|�M�i;�H��=(.`eϪ&A��9(%�3'Dz��f*��H$��}���\��%�����E�s�I(��<]�9 ;Լ���~�G�ݔn����wn�䣎���9tHy���pqXM���J�Oؓ5
*W��3�q��+�y5�+y�O�Cy�"���5��c��6@m	��N][��o^�_�HN�y���u2@�S��'�kU=���bS=�F���ٝ!N�Q�8��]��!JK#]D?Q)��i/�zJ��]�Y��CSeZ���^�n!���6��
{)k1U-e����_�����D�T�g��U��5��|�'ā�˗�ٔ�&�C����K�1:����ǔ,����SnV�p�A��H1/{��Ӊ�i��<��,'���Y=�>|詙����xO��U�v��*���Ȅ�hy���bn�&�Z$���<G��e�(˷u���LL��D�t��(����%���?��d�ѕ;���}��ŰƎ�v�2=צ]H�o Y<֡��nRk�l0T\P����t���L��cL5��Z�?���V<�G��))�@�����`���:�[$��S,y�N?rA4��s�A����r1�NzV#�@oxjT����к~��z�'�z�tBtyȅ���f+QU�i�+%Pf��<���o}#���Z��O�َF�Ʒg�L��Q��"\��?�W������1i�{02��i�9�9�('|f�3���P��ծ���rG�?��ǃ��/KJ$&3�k2��!�ք��᭒B�>���+�o��'MGB�����Wd�j�@�����}��4e�q���-��?�?=R-��U��F6��r8�m�&�.B|���.A�᠀���,���>E[��z���R^u\���̢2�a�ɡGh�0'!]R�3pe����.Ҟ�OW2n�}��A���-f��g>~5�הpӰ��uF���MR	��n���}��"ݺ�^�=���caN�A��2��s�%�����D�_���ʬT,lvC�I�na�e�Ȍ
c�Cf���]���BȈ�����'�~#��:��/������EpO�Vj>�~m�yaʁ���1��/�7h��#qkmI�`������x<�͔��(�A
cJT�-�ͺgV�G/�j���a�z�k����>�־����%�V�����(d;TW�����	�m��07���	+��+��Y3��ռ�y<̊���p�0g��A�U�v0i���Q͎�چSn>�u���v��V@c�,�ϳ��>{LT陃���pr"�վ���{������jH��M5gaJ9���}��=����.(*�/�v�[*���@:y��������u7�PA�Sa9|6W�I� �����������]����U��dǋ�7���G9�ӥJ�6g�3s�ܢWpa��O���� 0�%�L��\��mr���fVp���*؏�e6�hb|0�G�$�ñζUy��Je��'�kcT@͞�I����C��ӊ��47�f��������*Y��kw7��G��s�;��{�U���JH�����Ƌ5�z�;�_ο�������-������Z�Yn|�y�_��*�q;+ቃᩐ{���u>��L+�ܓݾ�����XtyR��ۼ�I T�vTۇdRղ�6���2�Lz�[h^c�_��k'���4k7�ޠ
|m�*�P=X�D8*y���
J���a[x��l��)����&�yd�He��ԍ���܅N��~�)�;]�a5�:)����o�7·v�~'��k�g)V��5�9�8[��������P���tz� �L,ʭ��|����}5�q��c>VO19���I=i��t��P�����fx��>�3�%gq�8�� �ԝ�ׂ����}=	˞ՁT�&�,�j-9i��v�n=�z�V�䔵I�Ν=q�������@�N�Kf@Y��Z���}qn��
I�����4���X
�m�~��ơa�Vg����6M.���=1 V0Uh�V����Cm����?�^�X�Y�VTd0���3�����K��|��Hz,yDH΃�Uy#���Ao�W�l���d9���
`�I��l�y	���9�r���M�Z�"�����26C��(���>��z�\�����LM��9����i4�7�
.}�\���I���:}�|�%�$�V�)� �C�Ҏ�T.Z��<� w��2h�;���3;X0��1�����o�}w��A%z#�Z�Lǝ6(Q,��0~��ak��+�$�J|w;x��BE��#?t����t�	�ž�����8y��Iث�*��R��1�;�p�Ia5��W�T�-�j��,s��?�G0�B�o�+�R�)(���ʣdp�iU��)/�4b+�ǲԌc���M��mJ=�>O��E��fD���c��ԩ�mR|�!�^�t
����L0��ԭ�`��'��L�Z�:���]ϩ��������p�������u�b�:*�m/6h��D��h��lJF���!֗eD[6� !Ficǉ}+�(��
JjGK�
�`B {[lI)g@\G��30I0�ܽB~/q�k��w�VYz��A)p�T����-�f�Y�<]�o�ƂG�\�p�N���tn!H���#S9����2h���T�5<�,�h1Ms��	�[D���G�J�Ʒ�ϰ^�e��Vp����s>��+��XrS?!�����|<�	i�$�Ն�{�}��8��:�ꫥ9EMy��VN�k�v������</X�4&9��U-tL�)�*��ܛ=� �vP�r����ش^%���[~s�k�� ��C{F�$+k���tZ�g�c̓��6佌YC��'�L�bT�%�O��i��35�
�"��Q#�8yԌ�}?ɏ} o\��G'���$q���]^kn�\���ڟ� yr�����o�+J9'����,�	���
�T�������"��7~~�R���~��/@�0�h�I�Ud���J��3���^mW�0t��8� z=�2�$�,��&0�+�{'� ���)�:,�ᮐ�5A3�я�q�ib2:Y̏�����,3��˅�'K_�EFJ�SW-o�#&.d�e�"�~&S��ݢ�֙a���� <!���"�QMN9EV��d��gK�2��n�Ȟê-����Q�}�	y9��\|i�J�)LG�J�V�;I����GV�N�S�H{�H�/o#2Z���Vla�B�����۰w��L�T����3��!2,;� ıT$vaY;M1�j��7�e7f��� `%�N���X>��žھ��d�I��fT3��;<��;��eaHe�9�Qfº&�Yo����c�aM�2�&��;�v&��������� D���P������\n@��"!o����'cUNs?�������_���|P�����Q�C_=$z}��Y�ר|X��rG��u���j�u�T�[$F�øx��UۏÍR@s *l��#X���r��e�p��y=�wu�].��1^���o~ۉ�dC]�aX�����-S�U����ܗ"Y��y�bډl$�տ�o��)}�r�c.���,<ɰ�k	�,����������/&�Y�C�w\�if�U�q$Ļ��N�k�����xn�dD����i�!G�4]�)��kT�y�q^[קMId�@��Y�B�i���l�� �1��L���t���lS�a*F��c@����Âֶ�^�El�=X��͘�1�f�#��<�&�+]SH{��xH�@����TgPcG�Q�,(E����l��Z��di0b\�ٳ
�x?�T�G�x%Y0d.�#i�}!�z_"��@Tw��93 �<��C�컇Vxj��(���Q�b���òQ6$����晾.�>}^��X��nc���Ďp�5�� r��T�W�]Ck�^�a�xaI����T�a�
�`�w9���ys3����͸��Ͱf�Am�]�Om&wh����~k�f/�wio��{�@9?����ҫP�Sd5��E�bM�<��P�$�L]���.3Š�3h*v�/�4R����]���I���m*� �_G����R���!6��	�i�L �d6����v����]m��^�qx0ycvy�C�>�x�zʤ���z�F��X�a�~���zM:_��OM����L'�Y��*��,��V�P�-�;���9����V2^p�F�)3�ڕ"[��+?�������f����W�`�w$�\�J�`��gD��̃>c#=9B&����c�ZX�Ղ�ug�&v�����:>�Z�p[��}U�\k�e�m2�yՓ����M;������3��J�K�XT�@��z�J���l�&��b������I�w�NȪ%Rg�1�*��~ ��!�% �����>�19n���W�*g1�����p:����)W��s>� @�a(̹G�m��k� ��
�T�����q`�t�n ��K��Z�x�~>�f�+֛���+G�ԁ��|B�\-"?��U|��v��QnvD��: �3�+�P��D$ƹ���@d��zjУ0�sP�@���%�8�D��,��gEr{�A�V�BYa:`~�:kMȃ)F��_Y��hP�������O��y���n8"/a��V'h���Hܾ��φ�И�Ut���o����H0X�,��A�9��Ӫ��׷2ٚ�=� �����z5J,�A��v�D��������֜hx.RjH˪��h�w;�n�Q�@�B}g��渿g��ar�B��3���B펇��/�� ��V۠!�ti��^X�+6�2
9��d��nR�� �1�UK�=�����H�m�K�"�@�{��0��ڲ��D
��/��t(�Netz�n�=U����.�hV�1aB�il\����o&�G�j'r#d���x��<裨�������
�CI�y>�΂�w�?�����Al1��N�Q��K�>١���Ka<Hp�q8�}Y�O��u���	J�bG��7a�;ͺ��g�o]�3`��ǘ٣W�3�=mK�w�aJ���F���w6�EP�pI�&:��]�#�bW�T�a�BO���f�D-]���z֜6�_rը��8����+�`����W	�����m������1*ҘDt���]�>k�y��f[E6��9���,-��π*a�6�)G���1�"8��7��t:��:'du���]�^�G��x/Kq��΄���&ϧ��҄oR�	&G���d��+ s����SQ��(�H�[&�@v��m��V>����um!��Ln9�w0k�+���Cc�e'���"��[�3�_�V�7fB�/���m�r�bN�����< ��L�[A�G|�+�4�
��tu�ʰ��HP���f�=�<�!�H��GŤn*:� �,%@_i@���O��b|�[��-w�u��[�bx���tB��Ɂ�6��X/:�`�G�kf��c6��ؽ������ʹ��K6Y9�<a+󖓖����FS	���KVY,��a17�;���p1= n� Wp6�\�AR=��c�'�[H<�Pz��p��Dc�j�9�u}��-J�} P�ڝ�?/����]����R9��3o���j�b��*?k����D��k@.�豬��}^�k�FN�`|,UtG_�Y���Q�}�뜦Y�_���%��EZ���D:��*纞�� OU�IM?�8��f\�ͫ{��{�, QK�n!]�C�@��U�.�b4��� ȭ�����$�ӄ�a7�ǿ���Ocm(��Ore?���)���41ǯ%ngW�YI����Q�O aG����y`����`7�b��Ÿ�;sdD��fo P��r@^��:ҿ(�u	Xn%. ���lYR��KU��.;DQW���}�r�<~���<��c�R�\4S���$Bq�&�&�w��\��5�zU�����y63O�jw��!�F����x�^=w�#'?Q'�u�8׵���b�r5���N�nw�\��H�:=�)WӀ���*���@�9�#�?ҡ��x4'o�_uPUBޯ��3mC98]�ᰨ���̢ Ld73,�Y��0�΋\fŕ����+0Ð��
X�X��]����\��p�Ƹ�XN�q8���ҫn��>��K��JXlxVHYEB    fa00    1e30%�Ȍ�%�o�z�K�|�`X�#Y_W���uzs5!�����'{S�(U�ݳ~��p'a?'��`�s7(��~�����tF��::-4e�T$㥳ɤ��#{�_��`����|�}��n��t3���'�J:�c��,GT���Q<%�����������~�2U[��'f$��"��S�-S4@�����&}m��i.�a�Q@�>:��F����v��T��Q4�$�x�p�jp�)��ټ�o�P������!��:�v�g,B�_�惏z	v���TA%�%�-z����.b�b���q��>� �l�U��6������^��bN#���Q���S��[9��	t)�����g��hm�ً�4��~t0���v�FTl1j�əV��I��!S{�-��R�5�^�I�y+��ꄩ�Q&��b�f�~�yukޒVik@XAa4�蕧";���w� %a�W-,��_2Y@��B+x����SA�|�QC����G���ae���>x�Y�J�w��پy+��<j#ֈ�!R���d(����uhOý���
)[[4h.��\sߴ�t|�{s�v�.Ʊ������J���<��Đ!�b�u�����*��OV��T$XᥙWt!ø�u�u�mJ�)Ca��c��KT��O��b�in���z��N�`�Q��^#��y�'BH�a�B�<�݊��t1������U��I�C]�ÛZ����H���K����:R��Uշ�K�z·|hB)�E�~�7?��a8\����v\��t��U���d՛�
��)Pal_i�4W�&'��A�vƓ��E*�Kr�,����w'�Y�ƪ�4�[�jQ;�bj�G�\vR���ժo 	��>����7�=䉂&s��K��YAB]Ǆ��(����[YБ�ruH�=�ލ�R�n9��k����+��(��� ��8�H��c$��,bb��W��TqGa}� �4E�r�r�NU��(�M`'��'�R;k��Q*:+���>�/T�boFE�C1[E��&뵕�{]"Ӕ�3���V�V��ܞ����GtIy��Ϛl�+���~2�57�,�={���	C�^��7��j�=�P�>ї����.ˆI��G��u��j��~ߎ�Isx�ٚ3����j�hl��#d6y�fI�07C������d�����='#���e׼-㷁��wI�b7T�c�fop���X!V��Y�ғkVKƥ�����w�eĈl�^��|�7��"@�X��ʍ4���?OWR@S�۰ɂ������	f��L��9"`�����g���XM����i�nS#O��{��{hL���%t��	P_��`���0�	_z�US�x�6r/'��ɽi
!-u��K�ю�.�ϐ3������Q�Z<��
6�2�I�b��6�žkPҬ������W/��3��f&��"�	TM>j���>�U�C�����ǽ^x��]��CY�^H��A��J��!�G��w7�pT����$/qܷ�]����J��'�w�p�̲|��x��ߤ�ϟ[_�t�k�`RH��N�X2��,�K�W}9�W�\�2y��fU�Q�ǰ���\k�s�m�e�+���
\d��l�zt/f*��jp��T���G,�<i��c5@��pW�����Aع��Dd��&�=(��}'��~��V����T�`U�k$~�o�͎ r��\��cj.�nr%j��-y5���J�3{2�!�Ӕ��e<�4��Q����Os^�����]n�̻����Cg� Q�;��B��������l�'<t?$�+C32�l�t��,,���ɗ�&b ����!�d�S�#�bs!�a<�/�e�2F�� (�������\��\`:���F����H�� ߜ��bD���V.T׉�Z
��׋�T7 ��j���ƫk-��uK�\1gƢg�\�p��~��K��b�Ж!Ʃ��,eƨ�Ģ@�L�}��t��占�2N.� B��}�1�-��쨕�0��mL�-q�T	���m�-�3pT*������I��o�M
�mV�{�>�F��`�������^�w�B�I�L ?pU��d,��Tn_�?"�I�WF���#I���0��;aׁ�e�G��YS8���η93���IV��L���4�Ϫ����an<E}���`y�RE�RO^T��������!�7{���E��O��ݠj���U&�Pm�b ��M�t�b$!x����`���a�;�P�G
fp�j����i:,4�.�D9���Ҳ���}��[8^k�h>jaU�!�uZ=��Ti����:����ܞ&ыXA`��x�2;�P�s��<x����U�J��- �)TFKH:�,N���X;�<�[Jin�g�eϊ� d�~�r �&�2}S��+^���Y�!K�D>6�(DQ��Ҿ���_׹͛a��>�U����]�y�,��5�i�V��F&U�V�x�*%�_b��缺�)��%��_��:����TI� aWO�j��\.��kB�>A���K�<�e�ң�~m���?���1�eZ�m��90�;0��a����9Q�^T,~l���$�@�_Q;s���<h�,ڃ$�"�nQ��?��(���nj&�?u���EJ7��|�ž�q���\ʘ�Mu������N%~-������Dr�EP���n�*`�۵[0���ß���������g'{��r�S�;lW�(�u��_�N4�ۭ�a�*�W`b܁m��H�P�v���	�T߅�V�ne@��2���^��ڣ3~����~eQ��FNި�c�u��o���b ����'����S��
..��/��=���/�h/<F����hXY1�=	������p�8(t�k��pU���,�5�(5Ro��`%�᱉���m�v�{�����< 2�I� 1�����`ia6M����Mt.���c�]��7�̞�cg��oF1���,EDSp��`���	��tV��=�	���xD���z��3��ک|*K�����{`^Z���L�-��c�tF|\�����?:\¿�K.):�*H(h�\?�?��qS8�@O�m7��������m���+�
F�zq%�Ό�Iulj���|�}x�&m�Ňܒ;�{��ڳXh�Y!1"(�Sʲ����_��p���c�.^�zS���<�P��ѹ l���i�ǇM�	/GXz��oՁ����g�$��˪ #V�q�K
:��Q5�H��{Mi:\�oo
�*�X��rs΅��'�x�u�i��V�Ģb��d��ʕ�x��pU��b{�R�R<���:���v�h)�b�_G<��'T_J�)�"M����"w��Ȇ*�׾SU������/����ӡ�e�E!��.�W9QZ��jg�0�t���j�� �4|�*�Z`>A%�)׫��@Ϥ�����i��?�|b?-]�oF�ջ����@7����>2I��͎�'/*���[u�3�.�%%Ϭ3��5�2>�I�3Z~^��vo��#��ZXb�خёh�GN_s�#�7K6�GMRp�����j�h�w���K�ñѝ]x&����kX���&A��̄�O����YK��Y�]�o5�z/C�t�"�
k�S�N��=����HdrK�Rʖ	�
��0;:�Cu�iyg	���c���8a�p���J�s�<͈HBU�yfٷ�Gj �+IG�ML����G6~H��~ؕ	M�߄��}9J��]������[Y�܂���U�ݙhdh�R�cHm̂�)��s`H����Ȋ
I�K��\\	^���.=_S���╟��*LҔ-ˑ�ikn�w�j���"�h�M�rNG01�A��S�T�1b�~I6��3�Po\U�GB���J5~��m���cO2@�����&�3sT�������u��K�J丞�/��|��f��ǁ��[6�y��I�P�+RI~P>��-hcX��E33�t���4 ��nVpm}~��{}�k�Yn.�	�A"�q�z0������ɵ�c�2)��
9
��ul[���8N��K��,|�u����[R�L����ˤ7�t*�n�N�dmM+F��#���%�R@b_�<J������\��%,HS��;����3TW�XW����]���X��c�#�XyS�[�X���U�,:����!��`��gMC��&	Z_g������Un��zj��sA��ဗ͟-� kiyGu�� j0{�3��p��
����7@�7j	�BU�u�s����j>Aƃl8�����")�D��{�w��&��j���|b����%�D2���ܞ̤?���O�a����.�~�d������κ���lO���1_�h����lH���5�ҟ�֓�C��~Y,��S:�ɥ���ty0�!�wq�Ŀp�
��U��8����dV�L����#�T�Z��OXF䆣:��4�"�L�_y�}���{��
�TW�ͳ������6��d��b:#�vD��Q���2G7Z-7%��d����z�,5b��b�gb�-n�{�f�ڠ�8D:�I��T�=�-�Ε:�?����q�C�'r�_gl�)����0\6��'����y�#p�����h�
q5H�T�{�L�[([-�M�����p�mvO��k(S��-��2n�hW�s�|J�Fp�dM��������2=�!�>	]��d�=uDR�	�(��8R7����.�_�:F܊Xgg�>�U
1!�^����Y1	D1h�g�'��U���{D��g��.	dl_!�m��0@)g���*!���*�s���y�&��Gl��WLG��z�z$��TxTۅ��t�]��s%"�2��ŉ�q��/�$
+�KT�0G0n1N�%h�;��P����L٠D��x�aY���8�we�`��楜 }����Eo<�'?���+��ohv�Z�~�OT��"G���p�6Ԏ��fvyW�[��l��c�_>I�&�m�z
W���w�%q���O�]/��E[�m-�ZC|2@l��o9�ss�ӏsCW����!�m�͕�����,>��^v�+%(d�v广��r���J�E!h�	�(�p����,�-��m�(�}֌� �*�Lt�f&T/4�E�P�7�Q~�-��ƛiR\���]q�Im���!�GC��/�G�w�g���Q�@�7,�,�0"}�u���;��!ϡT���i<�B�B�h�Ϊ���=�t�ogJNp �30�JFI~L��'���������^�H��H(�ȉ��<�v�:�AdBn�$fO�8-Sl Q�����l�޹C�r�M�$��>�!i�j�Ht�6�|�oڇ�ҀmH���� �Z�J�{_|m{�y:��^�T������8>^mӿFX���e��Ԇ���896������Y���2?/'��u��o�m����+�@����'�BhD_���5�k�|yo7��c y+��m�E��4���K�Uh(韻p��^�q�R�5=�w49�A�:�ea�ե��C�~j�F�Yu�eCˏB_���7w�-7�@%�.�v�*�%YΌL���o��~�1��t���b�h���E�y'�S�e���(����|��m�4�U>Mzb� v�	��4�Oi�G�nN��Ƒ���a��������_��=�'�X®~���X�7�VU���G����7.��[<a�Fe⇉62��C�Iö�Ɇ�*��$���3�}�;��
��3^TL���;e!�G���7�Y�O1�X׻Q,�U�M�<��*�o�	�t���t�Փ��O�_[�Һܷ7
�������	���X\Sr����'5��q�n���<{��mhҔ}��Z��l��:�5�ߐu>��㗧vv��a��H1���+���u���h�z�0(�&m.��A���h�6���}I�'N������c#�,d��J�U��������墓s@�\��nLh������K�����Z�[�#{	_�[�%�Zp2��@�xYW�5���ʸ��J�'�t�J���Sߓo���Qx��r�8���#�����Ey9�M�8�@�kʲ>J��{	�w�vf106(M�e�DiƑ�h�hM˽ᕸ �r�i�F��@���Ms�.u�%0�,�\mS^p^�&Ց=5��t�3@&-oo�C��.����o,����6�1�Q�W�Uԩ���ۼ\���@���i�6�%�W�]��x�p�+-A�w�Y�DbH�i�i�,|�"P[u��1��2zV��gSɀ��֯��c���u�h���F�=&T@� �B^�r1��q33mF�U�R�ޜI'~�d[����O����U�r� l�1��Ҧ7H�ʔy&7{�����w�|�9�� �-�;L�R5���4Y[�w��sR��5��Aĺ6�47��,h����_��H�#Jx\��Mfh�0ǹ-�M}�:��7S���0�S�23{��C9�ӴS���%���_�H�j�iϘ=�����s$��h�C����6p��*���Ғ�^&�Q$�\dR���ɖ�i�3��.P�oy<X�V�.���5,��^*���*��DP����gV'���<�]���U�&=&�G�'��B'��p(�MeWf��Y���>����T��	bzKߪFP�_ǂ��&���D��-�5��_K73���_��d�^S-K{+�ǖ)kI��l������t3;��uJ%�@�Q�ƈ��W�������g���,�] ���J�"x�l��I���rK��R�c�[�%82s��k9�Sk���DC�D���5�nj	/7�)p��9�ݶ�t�m'�%�}���
��5��
3�B��W��[�Z��4S�Q]��K<����5��y���8!	��6������]�FJ�q���)�����r_�X������6cq �{�C���?�\/��g��{+w�ԊSI�=�� ���(��ֻp��������w�@my��B�_�m���uR�װ)�-�լ��#���B�\0���b��Am�K�y՝!U@��7�bg��~�ï��1���B�oWٸ�
�%��g����*a�)P�`��F�k���K���}m<^���D�:yc��*%H�]��l΄�!|�g[��G������ML�����ź�ug�d��vYe�Px�`M(�H�k`�_���gqY�ɐ��<�J�W���OL�5t��Z0��W`���s�1Z�hP�dx��o"�G����?��n[��A�z>叿�kz�d�����U\�&B��3�Xw���� {�?�0�|�AZ�Ik���|T�'h���~v_K���D�6���8as�$�k\����s_OT�M��~���պ[ ͡a��#�T\O��t杊�>�����qܶKS���+�ظ�-~t�����|�D
�  �1ЎnO+���k���I� ďD���;r�%F�Y0�!5A�q�U��E�M�'�18�V��x�i�g1L%���
�EK�HB��5� �*~	w*_e�W�Ҙ e�J��
n���x�;CEV���'!fU.��I���x)��Y����V)<�uc�	��ߜ�Bܥ�Nku�v$b�W���S�*�O��\�� ���XXlxVHYEB    fa00    1d20�W�;&0ߕ����&�
����aF��~w�p�� 1�A�7�f��˷��!�B,gm@��DH��/����r�(���v�4��8lr�ti~©+��~/`�E��0(-v/��x7�'T(O�BW��.ԫo�W����>�BXZT���@Vrc���ܩ�$h���5*����Ht$��˕\4ަ^x-�N���B�4�'�E��d���N�Js�Cօ�By�>Ë�P�+�.���d��"o�Os��:���2���*%�Eo�aҴ�����>S�l�H��L�sV�)�2�n>/6/U�1=3�M)m��H=�P���T�Ð������J�-L)1
Ԃ�~�*�{��О�̷G��J��!F�uxYg�S2�|>�sK����^�QȘ��{��Q����<k(��NC��`�/��F��kS�,����od��-�vE|����o5��XiL�\ͬ[�5��?�E� o��Y8E��
�dp�'C9��w�~Ԍ�N�J�hy���I�<��3�*#��d�-w|�Rb��F���B�M�}9��woG��d�� &��X���P��2�H����u� �}�G1���a:��^c b�<ͽW��IW��u-�����d\�Df�P�g���ϼ�g��zp&�#�Q�Ą.���OC.㏈��ȹ-빯��H-&W������l��Vs�޼�,\r��0����C��w��Xy��5� ���lF�. 7�_��������fʅ�M�r�lP6F�lS����p���:?]ө���0c��Zyp�C�syұ�@@ �0�1{���a��F���Gt�w��9�t�wQ����\97����˧P�Q`�A��b`�KƦ�6��#B1�#����6�3�3��|�y�!oa�Mm�KBUa�]j	0� ��lץ���:��� ���(�Α
xd��o���L�9 ���<�eT��Õ�9*��sG���u:�i�42���ksPjh��.��+��C�M6�z8�1~oplt�8���Ȑ���v�n3T?���*^��@&|i���媝k��m�S�u�|j���񤷽���}M��<i�G�D�0������������� ~��@�ͼ~-pC1q�ut%/�-t�P`t�	ۥ�[:���Y��9b���A�KoeL����|��}f� ��6[	�?"t\�j�1E��G��$�"�F��}��J�t�J�*T��/�.u��7���/א�Ye�?�M�����4���G��-�ƙ���@�v�S�4���0�b���K)ۉ|i�/#�|/�s�'�:��t�V��a��!p�yA�z�����fsy��^�߽C���b2X�4�!\��;�H�����Q�5�Bᡰ���'�s��ո���
6��<���QR�N�^�Ag�ם�3F2�p���}rI�D/Pkǜ�B[0���1��
��_���U�4�+��x��ґg�!�tm��c�N�Xi��۬v2a���jn����c����m `��'{Y�Qs��<X�&�'��}f�Z�c)�*�#zn�w�7�rp�;8ǹ�EQ?���s�y��SǶqU@�	]��c���S�ƌ�U-Nk�,w J�澋����_@H��*"7-bٵ�� r:EN5f�dAR�F�Ou�"Vw�jC�m\c�}W�	��E�EDV6��H2L�b��Vw��>_�6�kHah��f�Q���(dF7���g�c]�f2��$��l=�5�D�Z�Q���,�>�̟�Gk��Y P�&az伾|��L�IK�gz����=��5��Fu��R�gCk{��9�� ^J������p�b�7<m����v���F���o՗v�������.TBD7��,���?�M�_�,K:��4�m��-L!s�[���	 �efE{L
8���~׶����m��U)�K�k�0�+���K��%���ޡxu�8:Kq+A$���<*/��&�w�*P�!��ؖzn��q��qM��(��Ɠ,�yR���boM}�;�6Z*�̟���J�c�uyɇ�5M5�0����Zmxm�#|����������8�{��lN7�GY�Su��}D���M��t̒�ZI��Eo�mĢ�Ȓ^H|��@V���| U�y��c=ˁ*]�d�@����[���ҿ(�gz4�z�}����x�UM�0#X��u�3���[k�`U���6�Da��ɝJɭ����Y��咬�O§%将˘���`���8d�s<9p$�y��I��!�EX���QW�F���o��ת�б[�}�P�.d�T�tw�ӗ{��P [�*H?d���q��blӭ���ɍ;����N�:H%⎻
��j���N��-݁����3��q��U��|`�O������g���WtZL�F��g�6�d;����-�;9��B:ӂ%b�.�vG҅�_ Z��>\ëfx�z*4߳).�'5�ꌈ�%��4�eoS��Zx�D�n0��}Ǖ��-�2o���2Y�GKbtآ~����t8�l���g�,~�u)l�%�6']����^�ڒN2y�����H�1�Av�3�,��wq�ց35߁���3�:�>~�/��&���N���@���\(i�۪qp�|<��g����P�������M^�`��~�9�s7t���!�����]?���� ���@2�	�B�Jժ�+��(t���u�Z5��X�d�����f���zL9�ҙƨ����.��8>A���nVΤ���si�;@����S�;4R�`b�*Z����!3"~�y�>���Xk���8��>�����	��kɌ:<u0�4A"ƄZу(!����n�s�+QH%���̼��hF"IZ�,�o��X7)��7�q 3�OXڀ�
�~����X�t~����{N��`*�� g�g�k�l!X���2z��c�r��	0>�ވ�a�è�;k�y��̷d֗.'��hw	�R=�:���h?��oRg�(�i�o�y����O�A�� 	i�+Z\�י1��N�_Q�&�Q��i�o�tЮ���G�)!��	o����W����8vT%�0�����wU�;p_����Y��K�^���)� l���'/���ɩ�\+/�=��&�V�ӉF��)��¬�Y�rA($��qH���+�w�R�0}h?vHٚ��+\h���P����En�+�3��Bp[���"��B����?����C@�Q��S�n��=�|��J��ǜ��\��V��z��_��³���e�`O6��Oߢ*X����}��d���ߊ;g���d�72��2�vI����Ol�x[Y��+�Z�M!�����o�7[�Y�p,&Ks�Erj��ט��� $$u��hs���>�Y��|��b���Q�ݧ�3)-�� 8�l;;� ���D0iD�Ӏ}�b��=|jF�����$��Dξʹm��x+��M�V!���N~���F#C^��7HY���A]1��ǔ����6��2��~d#�RX@�H,��q�e�yhlh���tV�G�u��.e��J��Q)�n�{��|�����0�b(�7�o�!�c���d���g���/���10��hX��|�m�8o�����d���<p�b1a� �Īp����\W>�1�&����Y�_F����Ԣ��i}�;n燀 ���b��4�S�S�[�蛦Z�%xQ��V	�B�N@K��v$d4�o���w(u��6�l�����Ng��d2"�7�P����7T�����}�u�r�@"6����F��D�#������g�c���h=m������f���dUz��ծ�<О�Ǆ�&����o�?4��$z�uū�f���U34g�ڙgc'��RR0��������̧Rh��$��d�����ImT��v����{�8p
�2�)���wѴΥ��gn�G�	���m���k��X�[��w��ۻ�=�G����k̙�����Z�2�M����u5�xD��nG�)z��E�^<���R��@J,��v*���TU�Ĕ9]*N�sa�fգqβ1��z�.��������ey֚�_j���eA�F3~20�Տ?GhZ��7����<՜�y�e�;��]�G�U�5�}�����s��������2�ф�����E����}��łf���+B(Y|,w"�� �4fc�Zh>N,�Z�!�r���Д��^;)�� XP�����f�>���"�U�ud�Ҧ��g_�i�hlI��V�f�g�9�N��'���9��Ô]-�	��!���k���n��6��;��,��(?Z���ᒫ[7�6Xs}$�y�4���)@��b g	&�W9W	�"�IW���~ێ�:�O0��/��BBg�R��?$��D�x:G����963T��� ߍ��ڪ?�(�K)�#Ӧ^�8��T��^����N$i�W"68�-��~%\\����.ju��[_'������TM� )��hs�J�Ҏ0��
�s�a&uC�*����y����9�L��VzһC������ޞ'yrL��J!�K��Ļ�׊�(]��R/TV�?+��-"�P#�Ў�O�M�B�T3*l�Lj��(�`:��2�����"e7m���������&J�݇x����� �g�	t���J�p� �\J�����?����%BN$-����O>ɠ�9B0�Īv7�:�@l�������_t�*�?��A�p�cB�_�8���~��3ٝ�p� �ڦu����?2W��g��^>"fײ�V_𱬯:K{ۀ+�g0���۪-��|��%�$��AVݟ����k/�޶&C7;�&2۞9X5ڽ��Nt@�m��}����h֩j���4�Y6��nZ�]4k�ɑ���Of��(��l���{�Ub�'�<����wp�: ���|���(��͍(8>�~�sk�ݓ��ݾ(�Y
�"3���?D!�H��\�.��"�D�r��d�G���,���;����6D9
rOל�sz˙�J_�0nC�9�{	�K�F���d�?"ؖpe����
������@@N��e�6���tr��oT%n\��EJ���|xi��\(�Q)�p�V�Gk��Fk"%�l��Vs>aͻ�Х���qY������ ����9��7�Êb�l	�����E�6�L�4�Y;���A}e�ك�f���W.� ��=�Sb�]���{�[�;ڥ�p(��|١��OLh]0�z�<�U�����ʣ�O���[����}�sY[��6.�ܬ`gg�p5��B/Z���FF�"����"ggGq��3I������N��ү
����l�c<�7�xx�̈Iϵ��O:mX_OK��`?A���rk� 	�a�(�����T�d�W�7]��R�8�_�ͫ��+ˮM���Kt��=\�\�������h�Im��W���\���>�LI��N�
�f=�G눶G��
wR~Z|WK�g���I�Q�@!J���F{ӊ��'���(�E�>V�S�=�W �S�=8 �<C*�y��s�
�`���N$��K�$���d�I����F�w*�����_�ă�g�M����1��`0����|�!��v��9hӬ�~������8)/�/�=Cm�&^�R9�@?g�J	��$I! 'Y��^רM������S�`�D�=� ��ʹh]�d�aI�\��֥k�tɹ�)�rd�ߝ�C��!UV���	��7��X��wr�����@� ���M���8.Y��9Ōpc����z�s;����L4H{v$��H^r�Y��+��.x�t:<����Qhq��ZT4�q��B��F3��/?mf�
�$Q< ��� �4Vb�>vˤvYǋ�ڢ��W�J�x�#W��}�1�^1/{�V��OR�г7о�GUJf�ב���Av9���@ek��
F�z��@t�M���+<p���YGg�[R�[��M�X��.[�ꤢ	�Nfr�G%�U�c���5�d��}$/��T�A���:�m
�6u�b(�^����ʱ�0t��R�����-� UD��xi�J�������)������
�����+���m�݉�lI�C��Sޡ˴<yʨ:��hWz8���S�?k���ƚR� �LXN��Х|Q���V��ֵ��p�A��k�3��˳��8UH�Y)���0��)�}� v{h=�'�����z�Y1Qi}�U����G���QF>[�	Y�6ԣe�d1c%>�Q�����&����z����ʦX~�#L������\^{?�¢X}+ޓd&r5�"9}JxR<�c��>��g�8���⚟L8�IRR��wW��Q�w%>�jDT��|^�� #мՑ~�R�^��$�{�HF��%+k�H���v� ľ�,�ݙi�	
�.F��1���Yl�&� ]��q�R�N���Q���s0�m|~)� �Y	Z�C�޾�h�2\Zn��rv�������@�<índ�I��w�.�����Um��n��ߥ//C������Q �����F�(W�r��8C9���>)x�����l�a�͝ԩ]��ӈ�t�B��\�i	c�yvT�`^O�!��K�'��� Y%ތS�yX�f�j���V��(Ԗ��񛷘�F_��0��C P>�۸+���qק'�h����p��D��*9B����3Oz/^�FHK�3q �sc��m��Z�\��1�V	<���ɨ^9�(-3$�>|}ӝȧ5	���&�_Ҝ,X��{B��w�kk����Ƌ��d)�k��ݳ6�_�R>��ŭ
��n��*�r��O�*��y���ƥ�;^�C2����ZU��Q�E<���DwͰ�� �ǂ��Rg����.)zQemz����C�U�iSL䦊��D(���n�>�V�:�������7T��T���{�ղ����� ��sc:P��H�VQ��?��U����P}C����_x��b�E���}7i8L�����C�̣�+iMg�Ҕz0þŜ��~�O?{� ګ��0w���"w-��+.�#�����y=����I\,���l:�%�לs`��G��z�Q�,�˴g�)۷r����t?2��*Eg%ݲ���e�g 7��C!< ���* �[�.���cO�s��#�PmWt��t�1���-�y��p�&O\�, ��NT��s�a|Q�� 	��q��E��|����>�Q�'`�����6������;�a��w�CY���ƍ�9�[z��H�%)O�Nm.�?��h�������mJ��>�A����c�Zi��Y#��V���c�ل��gɫ�;|~J)Ȭ@���6@��`Y�?�/��a�ud����XZ�@i7��$
��'wږ�4	��`(�����&OF/;��6��	ٟ�0�8�XlxVHYEB    fa00    1e20��##�oF���1ұ-�(���]z���-۟~~��LB�(W�p�Q���B����PЅ��C[�%#Lv�8\�O�=�t��]�1��~ͱM^U��_/*0X钣��9z��pg���JKW���k9qO�KDu��K�acB���9�����P*a�Ш�����(-lOQ��A�r���S����A��[�\̙'Y��	`+I�[�z.eq��y]�b� �<[�27��T�.Ӗ��$x��t��#BP��!(mԅI����*�T�#�z�Q8Ѳ�	���?�>���^�βX_8枫X7�9,G�}t�'a*�ʍ'2	���H���9���ġ� �*�������.1��ԕ̥�0u�I�O��b4��!=�o���
����s�f���~ ��ܟ��ږuSD!�w�i�?�!���⬰BӼ����'��9\L�R��l�͕�'�����.|z;��2�wG��g�L�
�$�u����W?CYp ��@^ ����Cۈ���d!7�9�+ojF��`w���gaG5<G��eW��Ҍ�;b���s ���Q	�yι ��~a睝1V����pESy�ϐq��`2|$D��Vz�3X����̤������l��!]�{��LÂ��v�/��]x��\=�d�M���%��C���!���r��I�ݎ��>:��졀K'�GH�t@��ǟ�+�}JK ѩ́"�N��v|���C\��1���qx]Y�w�o�:�|�h�4P�]ǁV�]\l��/�]0��)����5z�a�.�M�R%|�ٿg�C��U��i|�Gp�s�����f�?'"ķȥ��H�)��QBC��)�����~?�]� H��K�n7�gW�<�ɞ��~���@���T����ZB-*g_oP���؀j��f��\�'tt��l�:��i�p��u[����0��s��W�N,�g�[;��;Y���&��H�dw�*���V2�ݹ�e��b���M
�f�-E��ǇS�A���]���Y(������B�ˁ�w�	�U�9�z��Ř:s�� ���x
�v�DN=���,#�;�v�%mx�M�)T�)%�*�A%�l'�Q~�z )��/��
-�^N*��շ��I�B`�͌��|���)��K+xs�B�&\S����Q*�-��_��1��*�js�Z"����9M���6��;M4�Y��f;�L�5���" o��N�kx����&�p�4A�aE�L�6O���o�0�����F�'Ci��+1C�3ӠB����!�e�D��`�[�fO �+�H��Q��ڗS݄�������8�G�/P��b���.���@�{�;�3Cn������C/)|����<)�3�b���zF�G��9s'/oȩ��
1��Ĉ��������WUBB�XKwF}-2;ơyy�?�a�������tB�,��I�!|@s����8B�2
y� ��2��b0-�!��~�lR�����m�����8��E�Vܝ��Aໜ
�)�/��Ǥ�iO���-TO(��}��c9-� ��R.�k��~��>"v�D���+���tk�{D5��p�wT��:�G�|�yt�	����2�pT E[��p1�K8t���3)(h����rؤx����
w��2��D�)m"��8_] �G_�M:�,��u���/��a�$�B@�ԫ�Ki(MI��ѯ��5 ������V�!����_�t5j���"&�TO���%u�����0h9�a�)2��}�UA_�`_�^��Ao����G�1���L^r꾄Y�����(��[S���{�|=?�����g�>A��͗[`.@Ձg9�ʞ@���W��G�����vP���t3xu����O^b�i�ҦM�o}e]�6���W)v�h�\��^��Eyk�}�N�M�\K/?���epSk�N�&�Z���Ȋ�7O����%�%AW��Y��ā"�7��@i5�.@H�2J���<���)�؁��^i�ldwkް� �_@����]��J�fr�~9�aɒ�~�Ʋ$��Ḵ�Wj��C]�a�֙�^;A��zF3�.H.3ԯh<����O�91��^��Ȃ�옅�No��%�Z$�0�������U�.�u�D����q�yF}��7��Ϋ�1�e%S+&S���g�^=�`��M8����NI�[�C��h���9] ǖ֨'2���<I8<5�+l�,�P�om�4��̠�v,�d����^��F�^f�'μZM���vC��h��7HϐӍ7�p��RbӦ��&��t���e�ə���7{��澢��Ǘ#�ό��E���RG�#�@��do��]p��z�Kˮ���
؈C�Z�z#���"I��D�Q��m��L��@!�4۾�9����v�F>',��3��BE$�����9�6;+,��?�̕f��
+��.9L����MG$Y�����8i�/�[^�b�����i���z�Rf�=a�����%'�*���r�g(�H'���R��ymr�9Є���E�l\�!~�V��2��j�54��F�y7�0VrL�K)��{z^e�� �*�L�,϶��um����邱�%|!�5��0���vZ�!F��n���3�@�:�f��:�������d��I����H�c�݋���I�9�^��K�����O�#5,x �|=
Y�'��M�t?i�V����;MՑq�㻟��� ʙ�D��4� r�q����%�O<!��=](4��H�0}�i���rR�c��ܥn`;�����V��0��_�_�K�'�����h�"��>����/7@@�j�s� ~��5��2�В�%�������L�g�*�PG8���-�tm��D�2�T��B�@�I��J�5�W�ͩYc�|y��"u��W���������t"�A�h�B��)�NY�������'�4����0+��\�.�,����Ɓx�,ܚ��%� !��W�nH�Ǚ�M�zKW਋M�021#�|hH��6�����&���*���N���6�)�цb#I.�̞��pad`h�� i*'�b!�V���du7��0ћDg�(Q��3b�Na�"̓8����yN�R����+F�oc��]��bF�q�:a�3��ɥ�U��l(��r��SN���[�g�<0����}���!2��.Hu%�(��H�&��J��f�M�%�o:�!��>�>0�d"����_>��CǎX�g�<I�V7��I�U��U&pw�l�+�c6:��s�;�!��L����9N��ڒu���g�xb������ƣz���n��i}� FS\�t#ī�� &#�f���	�+�Y�+�	xO��a7D�J ��ݶ] �7v����d���EP[�O�`�>Y��}� $qw�\���9,Tc�Tco�"'k�i�Z�b�����߰��Q
��
�4=U;�[��t`8܆ @�#m�p�O���Ш�_w�/���h� ����4AHD�$�s'���89cl�X�O!� aV��5's�|g.�Dh�B��0}�b^ׇ�R&{v�3���?oh�S��<A˵Ǡ������Z~���7�_p���	E�a� eY�^��r�������w��h�^�j��k;^��L6�!���� \# ��?�x!��ňSn�ĝIV�C�)�+V���&GFj�����i�s{j�s�nX�RLP�$��H�7b��$���ޓl��E��$��cSy�X�<|ū�f�/y�T����y��.�+OIiI�-��i��y%#k����%�WQ{�p�#�L|S�u|Ut��Y�e�=W%-��r2����9i�6�3��,e�د�Z��D���PN{����0ڍu�J�K= ��"��c��}:�G�	;�?�Tc�2"�[�
4\�&'�"N#�n���Xr���l����,�,V�*P��]��#��1-G�f'��.rQ'X5"�;����՝W�8�AB|!��1��s�FK����ջ�I��!9�t�Q
�����V�Yb�0��R��@Q����8�"�wǌ�s�nխ�rwKx�*:��~�k�/J�d�6*췓����$���nP�x�rk�5q܄~T��7\�LP�ݟ��e�+,3�1{R�	]�(�g����Ɍ�U�f���k�ә^�ӭ_����Y�c�EN�Ȼ���do���� �|G���z��>��k��(dvS����lOBT!���r�[���7\�:��Qn� Tr��/2\O4�"�z%��_9�EN�c+�c��쓔r���+�]����R�cw��k�&�������9}�g���x�[��/JI�1��4n��x�C� �</���!8|�&��$��Ђ��a��a��n1����s�����<���)�Ȩ�(��O�Jn���7��|H0; �R�|�R���؃�#���� �_5Z8�� Y��E
=�s�j�! �0�:��ߝ�����-�C����k9O� #7�Ȃ�lrW�~�=H(Ll` �
I�Z��=�+z4o�|�����Iɛ������X�L����x!Ư��?*��7��C}��|u8r�V� �qۅ����g�$h���G�萸,���ps/W,���Ơ��������c�ޑ{�=ߚ�50���5�}0x����9	C�i�ء�H�c�, v"��h�{ۉ{��գԄ/���2�2��Nl˰qp��|�s0��0I�BkQ��Ru���"r��*���|i�U'����r3,%&��C����i��[�h�@��cu�����$.��?���t�Ţ��$��g��=E�����y�v�ըQ�%ϵ�L� 8�Ǳڜ#,�<
�;�)AH���1U�.�-��r��Ұ�քD�; �_v�<�V֥hk_�,��Ձ�}[�yj.K�l���H{�č��.\E�"��z,�n�E�}�Tg9��������v{|n��%���F#i��p��ݔ�d=���X�C��x���+�=X:����ҍ��K��^��4�+��*[���Qߍpk0����P�T尅,��k�IΟ�Q"l�"�=���a��φ��-x��ڶ
Ȳ@֗%��-E�!on�lN~�g��2x9��a��H��nǱZ� W��(Q^�V���"�=o�9�C	���/�W��n{ �Z	����*�>Qw!�p�n'�;�ӝ� o�0�M�z�zh9�(��6���"
��� �P���1˴�Ѧ�
Ez9��n���-K�	4�J�j*��?tz�����Ln�%�W����$eI�K5:�Y\@o�'��
q�����l.��"��Nl��w!�%S��ҷ}f~�Y[+u���?N�fR�B&>�t��o���N��3�)�ig��{��U5�;� ��~'��e���8�}�?�]V�b
$	�j�W�]��__ى�e, ��f�g��$��"��%��[��bo�(�u�|h5�U�_a;�E䡋g�䎨u²4Gx�I���{���#��}��������ф�����O��dO��t���D�3�� ��L�-�B`~ R��8�������2Oi��`�Ħ����,�&Eo1D���T��?:Wkc�8�7 ��{�	����a{+1�7�)%�\OM��#�Kj��S&�Nf���9�y].i2#���{
@zO��Jǚ���ud��b��s[@��~�N˨�\u�J�s�Tၳ���7�1�4��˙���#�k��g\-��yݕ� �F���7��o#�]V�� ;����8iW�M/?n.����x���O�wG򸍷�Pa����W*��#��Α�O�Uu�V����8Ӈ"�>�����00<��%K��GY��8�s�E��
�T��A�^ʖ�R���)j,%R^Z��'�W�&��������>�F�Nh�jH#]����UO���h���=۴\��Srr�?���rC����z��E�5�W�14����%5'�_l��ړ�����k�֚)DU�׮gt:/I� <F���$#C 9��b�J�oȨa��
l!���eC���5
�)1���*�����r>L<7��}�7E7")�	�9�5XMQ�U�]��� �7� H�K=Oh��X�t�w�&a+���/��i�]��+���6s�<rc��W��.N��g����8�����L�q�aH}y7��|c=����Q�����ݣ������K������1���y}N�3HUK(lG����3�Z�>g��ڹV���.d��U�21]�f��EP���Z��%�\�b7l�{ZO/��DI���SJ�^\��`BF�F.a��\�3�����-�ukR+��Yr�II����fK�0��ԥ~�[����1�&�f�]4I�n%*l:`e@#�~��=�G{�U���7�HI������f�vV#��<N�L�q�n8��T.s1H�d[Gj���T�鱼=���pPT���W30�E
�+@���C__���iY����:�* �"��-�ˑ^EwM�+��;W�r�����2탖��d{֠�C&pF�F����H|�T������	�D�����D4�v��v��@��p�`' 5Se,�߆�3�h�!�4�M��z����#��H��h�V�ߺ�����4SB6ZIX��mLib$�������l,aM�3�OMX��
��k�HR�B�_A�R����@�G��[��Z6��S_&�t̰��D�6���-�e�X���U)</s��4_Mi���9���}����x��`���������$�D��>��9���^%�$x9�NӘ��԰/QX��ӕW�:�R���g�]�4���ڜvK�\Z�X�n~����ǰ�+�\I`#�?ǜ��r�%L1����w�8��@�J����j��儽P��#m&u}�$��S1����R��H�N�����9�	3��-0�)w;HC����i8ӿ�7�g!��2'�O}/�EczN�>R
�B���C:�4JF�����Ri����0�W��Z{�E�f˓Ĩ��֝�F�*^�T�(aA�}�ELC��~��,���s�jܻ^�������Dd�[�����Ԏv#�
L����5z`ĥu�`2�g3�I�R�u��h�ԡ�x{�/#�R�x�55�L�����'Zd�u�@<R��ה�a�
�r=�ly�!���3p|ȵ��㵸�����a�7\Z[C�B�d�Ӟ�5�\��prk����`�5l�X]�ŀ}�	B�ġ���fG��9���s�o(ǎ]pA���pv�����Y  �үAplg�7֢�W�+��)�^A-�;�m!c������o�� ʒ㼀���VKc�]8�'5*`;�vI����N�=P*� Q�ؘNL�X+�v�w#�E�obq�tZ�nbD����5|v竾�Q����M`!¶&�E�Zs[Á��O�S�&֙������B�Gm�S{W�T-󑋥	7Ő���&�S�v�g�_#w'���gHL>1%�����R
�ST�(Ѝ�X�"d����o����/�Y���Y`��N�������iJ��z(u�Ι�΂��&�m���4ց�\Iu�c<0/�����㙷w#͒�Wσ.�oP��ऴhȦyz2�c>H%��
k�oXlxVHYEB    fa00    1e50Kj��/�6��J���P�$�� �Uh�ĘnM�LB�+j�u$
�c#\3Q�vЊ�r����
��"�,�[3�6r�3!�R^[)1:���Q��Ro�=B�~����1�aɠC���/���^/��H.���5�g{�?�m�UZ��KJhd�_8, sV%���m�1A�J�җ �'ԥ]�5I�ß�_Iء�k�^����h��$��
.����ZE�~a[��~��O�' �\S�ˁx�(z��7Q*��:{2�ޚaU�;��&��$��*�8����u�`�
�F�Z�H�mx��k�_0?<~W�vJ5���.��,k>ײ�d���)��K_Cl�|&�R�t�>}�kR�+���ym��S���"�fGC�Ĕ��V�0�U��IH��LC'�p����h����~y�W�ӆ���EYݤ,q�����M��(7)!Lg��Y�����D>�b �W�|ny��\=|W�L�(� ��  7�I�%j��
���{���7�4uhlR}G�Y3[�����0Bx�<[Yןk5v�R���EWp��pG�%���F[��Ć�'U�g��;��ؠ�Z�A��ȕ�x.U)	�%qbꆠWT/�m���	�Nm�F���)V7��֍.���� �G�7��ΐ_��)��t��j�8��&z.߱@t����`�)��nՈU�}�O|���I  
$�&
Z�єߍ��w�q�3�BN�n�Ax�r�"z�0cq�w��\�$����	�tZu�Eu�q����g7yHѷ��;��"g�a����x-,��Y�N�qϏ�nݘ�7{��쉪�����?w��Y�NcC�Ѭ/�$��m�N�`��H��`Q���H�����I�û�J���c�ǐ����H��u���g#�|�ڇ V��*�� ��/�d��n�o�~E(+C/����h�p]�����)������d��{����4 �(�|*�����|CnS��2ZK'.r��]��&���_���vZVCX�Ia�A�L����q'�@��"�	���Cp���rLUd�6���6�C[&���d��0C""���d&s���n)=8��;p��f�Z�[�{��oZw��1C.hA��;��3�I��������U��R��y�n,��UxW�3Nc&�RFW
�b|� ������fTd��6Rx��7���z�?>���ˇI�h��2-�����k�O��/ @P���׶NE�O�$ �e�>칧@bI-Hɣײǩ�7���F����1���$5|~�+��|p��nfMS��xs&?�P�MX�"�I��[Y���6Cˌԥ��ɥ3��CśP�〪�@'�,�ȹϖ= ��fc�p�f��hx)���~���c�)]����l1(Ǿ��#����=L��B��|��]n֜Ď�&��[��]�i�欏ɲ����Wo�Y���x�1�PI3,�4�1y,L>�n>��x�ȸrJW���6���=�t�K����џ�6)�K�ѶD��\Ե�=�l�j�2�o������{8��G� �nf�SP�^��B+�����=�)^����Ȩ?0o'^��	�
@���}~\hߞIM3�1�]�e?U�XН�)}
$ 0�2x3M˸7�[��"����9*��ƉXD��G�o�X�E��8d�[�韋��[�Y��(iQ ��3���3��w��VY�g���hls�L�������AR0��u���W$)zN��M��K�8	�[\Jumvp�m���Q��8�P���F��x� ���&�#�u�E����-Ȕ5�K�3l��Ak��J8�Z�^����o���x�)'I�������{�jD4MA�^$�,�;I�촫��F�D��r'�n�ܐk.�	:uIV�'bEN}#�ݯ�lsV��	��b�R4�UU��E��l�p�����$�,�dZ��{�yR��E���i����Nn5�֡�(J�9\;旬xK� S�nN���H}�ɑ�M�J����c�B&=�Φ�'�����]��K�iZcz���_}[�˴rI�4sv#+.;fadĉy���*:�yI�Y��B����n�;1���"�D�mQ�\����sХ$�ϵWݠ	f_u):d<��﵃�3�O���3���g���4�7�ຠ�m8w��D�H��rZ��?�2�?ǹW��1k����fj1�|x��pđՓ�c�&9JuktނY�-7Kg���m���s�{�$N]�ߧ���ђ�"���6��߅h� �W#e��������RDf�.�
���I�;8�;�AH��U1�-G����c�b|T��M����,ъ9��`1����r��?!��e���CI<�̀_a���F�a��TћT�0R�X<cV:��V��E�
Q^��4�S�@I�ɿΧ�r�W������מ���LT,���(&N��5�7-k��£g�+L8l�jk�+ �������R�����V��R�`1AX&�.%�l6C�����gy����$¾�3e�[����h+���u�����a,/恅�V��)��rP^ӄ��xh�+�A@J��i��r��O
l'�B��[�ϭtr[��J�{����e�bD�{��`$^���#$z��X�����j�+ۨL��=U��ퟹ�҂��;�I��R�=���U�E�ݗ>J���)o(�~'n֗�݇LzI��i��*f�GB�v(�J��~z�:��kqh��lj骷�"�-�1��j�Fπ�����)s�)o�#��O��ԝ�H�m�7�H���I���wP(�W��n��$s�<�����"�ѧm�`�I���țkf(KG�h�#�x>�I�6X�JS:�}6����������*�΍��(�i�n�6�����e�m���No��X��"�����B���)�`eMY�FKs�*�����oF�bG����_ψ��N�`m/��w!�$���^��|US���&hmT����W6B>�h��4&h{��<�����> ���Ǭ�Ϛy���h�{�;�,C�+�,nu�r���r%���w�<�EQw̪r�0^UG�h��M2��V&�P���-�*@|���h������L�׽R�F�*�sT�7�v�_>Q��h����+�k�w	:*�";���͋nԂ(^�Zm����0���v���
�lY���\#
AX�?2��y�_xelɍL�:Nuu΃F�W�j�x�d�IK�����r`�6�lб1]\�kG?K<�750��vI��\\h�:$�FC��~��8)���\a�-�]Ô�"IO�����D .�S,"�1�כ�ϫ"n�LO�b7'��e��išT���% H��KOqHD.Y�_�8Y�O�ϜU9�G���f�-�ЍDP��8�9�������{^^k�A���P�Y�.7 �g���3ʹ�;��9�{g�ᕑ�IC�\�뫟�<���ؐ�%�3XU�Ov���\\a+tK��U�_���5�ʤ��<2 ���r<p�gkFѪ�n��q��jTG��\O�T2�����|O۽��,��b�.�H�G���Ԑ����()���ޓ�0�'�'����8fg��w���J�j��v?h�qGoR�,̶C��/����8���c��c�lR��+�|��x4� �Ee��BN���2�|J\|q����Y��j,����7��Yn��q@��#�+��� L0��U(��-����Y�3��j���2������L�/�H�y|ӱ�Q�Lzi��W���dl��∘f����&n�R�i�[��1�e_��΅�ñ<���򡨞�9��'AEȃ��.�����.���Ջ���ۘ���'�-�wm?�H�!���EC��_/\�c�."ʗ���u��_�Y<�fJ)����������k�e��$�������<��:������ �
�T^Ė̵���`�t�����d�T�ԝ�#��{2g_S���-Z8�y�-oL�dLx�z��没�C��Io�Z�r�nCv��J>�驸(��w�4`E����ŏ�VF���$hP�w�\������1�e~�;��p=��Mť��/�U��!F�)~
����?�9�J����\�N��0�ZhA��>��0��a���^hN�]B�9�w7���>$�ւ���[9���|i}L�
��r�#�C����w��:�2^b�f��mu�T(��%���� �z�}b=Бs�v��k��2��/A� B�M������1����t�G�ZSb�/�^]�zS�g�O�1MĹ�B\��f�ɞH�Bަ���oO��v��� R;I�||�9��hW��S�����_;�� ��!�v|��i?�*7,�B>�f�'���xwl���.�V~�>���S��/�bKm�ѵ�m�(gJ//P�k��M��EuY�����ӥtH.�P�y��눔��W���Z�3�bvD���2ĴS�Z_�7�]?�b�a����A<K�obΜ�Y�KA�TF��u9��"�p���
��o��H��]�����[v�R�7� �HB�I�َ�xw�w�0��B���);���WS*�8��)О�k����5Ѥ���]�����Ud��|�ͼ�+��H��=�� ��$��?x�B����!<?@\8V��=7�)k�'���`\�J/h�"�uڵ�K걙�y��D�����qtn����,Yx���ݻ�q�ݖܨs�P
��YeaY(�*"k]�Ҵ��X)������v��%9�%��K:MW���a&�QUB�M7o�Ŀ0N dҒ{������^\�Q��R.lp@~R���{�B�[�=Q)-�I�W�=):}Y�u�u�X=��'���D�i��1�M=�	��]9>$�jQ���d���;�ۛ6�e�@}�.Wg�_���&Yd�@�|�C��wDՋ!w�x�����މf�/H
(}1��R1F-��.�!�����A�j��F��W����XI�h���Kd�����_<����#Km����v����E���er
}���֟:K�<�J�鯶�X�nT���)���3���+y����v��HY�ὲ��w0��3�r��>�%%�����S���:r��><�%�������1���2мS@�9ϧ'��S}`��mA�A����a�!:����x�	t `���V��K
��1p��\U�;���u����1��O>��M����yC�n�Ҵ����tcRL@�0�>��'�[	�4�C.��+�� 
V`/S���A�kjj[�%�w�D�������!e��R΄q]���
�7��H�o����ϳ�U�ڬ�kN����[��k����c�9ÔzA�Z�j'���0�l'~�$��}���={������p_sZ��ì`��Dr����V�8���ďN����۵�D��3m��Z�#Xe+- kGn����é8�_���ᅗI� a����r�;�|���:M^iܾX��,t��ƅjZp���/�N7,e�UM��H�0�Ұ�c	�v�/�`�Z������\�':5[�<�n�ӟ���-��:^"<v��ߗ� o�Icj�%k�L|'���T���Ǘ��cn��}0�d�&�KՆq��.�yh0��Ԩ���wBE��y��Lv�]�����y.�f��\�W��kOg�GE��Ñ��WCMn��}ŋ+��+>O��
��y4t(�/��������r�����얌�Đ�P���3�Xz���ƃLbTinq3�֯$Bfx�&�@�̹C�uM3~�[eݯm���^'�O=05� �<�TXO;vJѝEk2Y[�{��i��E\���)b4c�,�q)�~*ly�_!YN��X�e��c)��e$o>���`�*T���Q,n�ur���m�����~N��c��4d&"T��ҋ�^ަ^SM�'Y*	��p����F�`��)�k\p���ϥ��o��`|Q|OP(��8Rw����3N��6)l*_,�H��ǜa�|H7��Rǳ�I#˚`�w���q�d����#������Q���9��I�i�9P�8�K�&x��H4�� (矏�ڐ9��P6�-uP�G���NH�S�+n7�)D�h��B�G]O�����V0�YK�H�#���-)� ��i��[^���I�F5H��-M�Y�zƔ�0'�,�<8���&���B6咹<-Q��$O���5V�dT�2����0����D�U�6��L�� �Zο�T_�=��X��Um;�f��5���`���D�̫��H�$���]YF<ͺ!��I �VO.=��Pnk=�9p��m[��%�Wnǀ$�������]��JǊ)t�z���jѹO��RO����ǰA��FeGA��K�sdp_�y̟2�/a�J�۰h�������ݓL3����"�ƃ\~�	}kr�q���f��՟e�b�pΉ+�'�8^�TU��_�U\�}����w�	Å(�@�qOb���g�sU딚��Q�	')��2NMy:�iz�ԯQ�ޜjk�c���C'�NTHP���u�(MX�*8��pؔP�����p#�ht,D�M�+Y<�V/����o�L��X�)���|J�
��=��鸎�D��Ǯ����)u��j�S��hVE��5ſ��7��+��;]ip���&nL[m8=�ܺ�nB�C�HH�خ�0�%���0��i�z:	��'����@]E���nUP}S�!�NRo��Fےn����Gҷ�d^f*��_j#U�g�^[Z�u=0/+��(`�n���;�>F���� E=�u ����$���XU�;�ޙvb*�����+�rl×
�|��HQ}i�Jv� ,��R�ȊaJ�xwM��Lf�9�U�1�,����M�D��,EH:�DSѩ/����ct"��@�sʴ]����׭�����!*o�è��m�G�|��!\Y�
N�������S��5���=Ꮡݭ��0{�Tz����2(5#��!'�X�l<�x�;�Q���4�=@E����T�i�L(�i�s_��������"l��է�#TB�x�Gr�5�<���j0����jiD����y���:Y����&jF�kl�~���Ʌ7�#� �I����/E=�`��1�o�ZB�/,��(5��ru�ds�����¼��ߴJ|�����@TWLFa���œ��R)U�l�����8�IO�@\����#��%*,�̞���I�V��	Yq9�Ȝr��51� ��vo #��H��:@=�G�0�9��կS�T����(�c0z�qsS��4^�k�.I����a��̸n� �R��̜�Z{�U��N��et�2m~]�Ki�U��.��YB30Ѕ���O�^/�9u;�%?�ظ��0���`�x3n����լ:�Jm��M:eJ�+x��Y7I5�6G���J��!e2q��,>+w>뜑oېt�YQ4�������@��B�:�N����HT�.2����Wz���VwQk# ���oO���L��K=��$��ڞ`�&���y���\�@@�삀,&'�ZN�53�����7��S�X뺎�#��_�B��+r�.���U R�f5߁^�si1d�y<����i"�xk� ���jT=f$z<ڣ�s���8�+�DM��J�VR��B ��|!���y�k��A��[�#� �XlxVHYEB    fa00    1da0�v�����A��iF�Q�x�U��J���M�\V��P<Sz>���<��&uz�Q����/T�K�2dg5 ��:
6M;�9O�Џ�Z�m����6''j�����M���&F8�c&Jn�\2g��`�@�R,��
�����PXϛsG�K���+�+o���L\�T�-� 	Ωv�C���f�X2���0��m��cX�-�C����ZS�`*x��0[�M.֥7I��c��1�ǀ%Fs��#�����6��4
0�� >��ul�+/��y'����:d[��=S��A);�U|�[�h1��bf���X=a{��ꁊ�w�����l�)y�*���MV��#�@�<�y�Nև�~h�6����j���L��ï�,��6��N���w�7�8C�H��s8؛���z�t��!%u�<��wY�+���m>�U���KC%���LK�҅��U����r?�[�N�y#��Fv�i�ޅ��^x���f״+_��t��i�zM��ɗ����	�����r�B�mK�+��e.���F����@T$�|��Դ���I�����	�)�{*l�t�:#̛m�m~鲊�"�*@��%�o��Ly�𴳔.DNȾ�U&�W��T���$�X�0�[΂�9��r�����CAB?̯,�3A���������ϻ�^��T
��1�-�B��zLDR#��*|N��6�ns�%��(:�9n�X�lH�NP����>�Ҩ�7�'���ym���ʻ�N��W,�we�&@��"�t�X�ԕ��7xOV����V�x�1�"H�g٬<��=�b�S�4�8��J�@��_�c�a��(.�qG[��c�4ߕ����IR����:g�U��łY��2�`CU�!��l������{�^Y����9��#5�������8vlZͮ��(~�V��8��X�����O<9��,���Q����ʐ`���o\��[��:� ���)K��/ΈoGO�/k%N�W� ��g��aڡ�,d^(�#rTz,K�ԥq�^�U)��U8dz�Z5��c�� ���ʴ�d�.�0&9%�\��W����o1b8�&{S��)Kb�袰�_���\��w��VAĵ߯2��n�XvN���]�s�?��5�im�T6�Kj�/�1�z�����		�f�H+N�e,�m$	$�|�x�Uk`▬��*�W-�濧�F�;a��4�\m���JQo�s�����O$��>�Tnp��d�f�TYxxg�ق2p9���^Qo?�(r#���}3�q�����m�-]���{���5��0�����Am��4]1�|�Y��`�����g~MY䗃d��Lj ���i)fn(y�� FW 罷pX�%�
/��׮8/� ��}F���$��_�3�ι{R�u�\oF�f�n*Q[3K>
�|̱��	f��R�����%A�L ��5��O�H1�l������pV�@N+��~_�� �)���2�~�+I���F/��o��J�.r4ݹP�P�~�#��n>l��p���e��S��R軮(M��Dq�U&�������K'�P'�u�����9�-�Uu�5xt��������5X�վ?ۍeΜ^��)��xC�W��0���'t���@*gq-?h�V��b���Sx����:r�RË�V񙇧'��d,2�#�$oS�)A4h�����}�0�7Y�}P@��i����T���/(�d�袲��-h��fA����}��?e~��ٻ��2�q�s����[[��0���E ���Mt�s�A'1>�S��u�~��z��η�l~%l��y�Sxj}`��'�]��!�͖{��Twe�?m��S+:��|�ϊ~���w��Pz��U�6��8Vq�PB$D����Lv��c�(}߱ �����I��k}&D�-$|��H�b�y��9A�������q8�����d�,$$=�&���m�i(���]J]�
6ާl���H8=]N��5�C0���4��7����,g�;v3�2O�ٝ�x~6g��f{f�>���Uh��M�=-(���5�J���+7��4�C�+�|��"=_��g��Uݐ�k�U����J�d�Q�s.���T�
E��;���#�:�����U��2W�'���aq(����Â��k�lt�!ld�ct`f	�h��Ԩ\@����w]�B��<��Q��#(}Ё
jHy�@�٥�����R��!���C�!p��)�8�E�v��T��R<��Z~��37�o�W�I�'��*���8T���e���R�2�ϡ����kS/Q�m��	���}镈!����$o� 5�l0FZ���d����Zپ�$�m���n�z���%�~���f�^�� ̈́#�O�i�2{4�Kn�U���,�j�/z/xS��xs�x�
�H�'�+>HG/��:��:b�!!��2�ޫ��7O�;'�j�坡c}3'�q8#ᓂg.4��Rx�߹&�߾S�Do^����Z1�3w��?$K�f�!���2-Ӻ��)2i8�=Ůt9�hf�SdЯF�I��wׄ�vCl��)��{o��I�h�e�c �z���Vc�a��#��.����+4��_n0��3�޷�(������@�yβ�dų(���
W���$n:�U�?[@0�v���6^^�s&mۄDa8~��l$�k�8��i�W-[{���Pg}�Cu���~n;�L3��Ϙ&?\:ܽ���;)c�Q����<n;�U�[ f�b`�����E�p�T�䌆�TPy6�eo<q2L��M���IV.čLM�:'�KQl�kЩOS�79ز��8�8��/�����|,� �ʲ�Z�Q�dL}^��:|5��ݠ*&�N�;9o%�U�\T���f�_���c5�
�%����I'f 2[�a�L/�^��ܵU�gc����c��h�e���\DR.S��_8�Ĳ�����O�Ҝ�&��gx��@"�R,�#j� ]s�4F}W0��,��W�#Rz�5[���O���"�xd���y�� ��8����>d�J-��G�A'���;�+���;�����Nje� \�\G���O4�*)���7�0Ď���(��I�H2�sʿ�&�|G� ��
���ėŰ�GJ��' ׻��;*�N���fw-��*��1�rvtS�V�s�a��I$�O�f?��K�s�6Ȧ��7��TƮ��(�D3O�\��P	LP��&6^�w8I+*^�م�-�M��V��v�2�V~���s����iD��;9�d�dh#��,,���3�Gq��^�T%:MƷ�O��k�)7�g�SV�����w�{{��4Q�Λ>)4���#���"�歇�?����Ce8�f�Ȏ�����R�ntxi`���˂�=x ᐘ�)��^��KX����	�2a۳��󱈰B�[�{9=x��Ac�ؓ^x7wg��_K��(4s_�1�kLbr-g1���h���}Zv�tb���${��°�}X��<0�5aoё��-�]���l}�r�������z΁�~��s���6rF�UVxjzg-X�dŻ�I��=v׳�˝wB
�|܏�f�N�dHֵ��xc�3R��$�cם�۬-��b�=1׭(U����<{�	��V_�#�>:�E��{����ܸ���i"�N���ͷfj��Tk��Rf��uY����=�����~ q������p-�P_��0UA�RT��m��p�Z꿄�e�������q=%0���k�8X����c��W4���������LKe�s���`�$j�\I�5TѸ�B���P�{+�z�ֵu� �(���Ν��	�Bq�����n`�9=�$���h�O�T��S+i��v�uJ1z`���u�~m�EP�VnG�k�ga��B]��t����n��]Tsp��aX���Q�'��-��"���o7`G�J���ud^�CH�ft�~�j^�nJ�&)@d��������ǐ&cc�B�v��@�Vz"0{'C�p�C�]������Y��� ����J��9k��ICiDV�6��� �\$��Fa����=;Ms�����c�b;�D�/9����Kt�:J1��Q�Jk�Q���c�W���<14ZH���l}Q�2Վ� �C�°�M�U-�}T�b��"��'.�ç�K^B�(����DM�IX�'! ��֐���t,-ެϞM:�eC*�W/8���_��]��4!b�9L_*~a�wκ7 
�UC�Y��no:?z(#z�0�@
��5�##�"���g�0���q���J�/h��F�c�n��\=�:��PIm��To�xk�d^�75�L@;�7�R��k��!'��I���X�%�$�#M: �$��4;,��¤I�����| {Յz�u���x�]�ވ��9�k0U�Tn_��p.L��w�3���H`)�<)��C������S�B����*�aoY�[RDb���������`R,|��چ��ˢژ����y �:�h�mA�#,{ޤi�A�ڵl��p��鬽IڵCs�kd��Jp��Q`禵[��	�����I�¸� Ұ�q6T Qp��r�������z����d���~ǭ��ɋ�q�(To��ӟЌ���.��l�bG�3���\�G4�w��x%Z'{{����fr�[�����|�t�䄬�P�y��YB��h��^��k�YzY�c�㱇�a���r��Y�!��>�gnoDBƄ1M�\y�X'��EԼ��H�����
��)��u��=6�F��{;����1;$+����^W���������(R2��/��ڝ�|-h�ovP�܃��zbS�5u ��N�n�k,�z�Q�gh��A����y�|����o�ې�ɿ��HB��m�3uđ�t�f���AZ�,b�o$[]�1�.�+P^ܲ����f�WUΆԵ'#�7S�(J =��s������[�m$�^�"�`��]4�nev����R�;�`�E���x l����"�H�rT�H�޺�@�d�y�n7�^�h���'O���ʊȾ�۠4l�@��9\Oh!z��$�I�!�)�*�`�!�5nQ�4h���nC��c���ܷk����w"p�;�ː*��_Sg_f�X�/Op�G:2������`��ۢ]�}{FȲ��B����r9K�R�_?md������g����]�8��Zd`�{��sU��3lUСi�i�j��*�F�唖���p<�L�g*խ�K�y��s	�u�e�M��1�1����r�Z�u�p5��*X�8����,��-���#���^4�%-����Gbx�JX�\C��쩸������vD����&S�+�^��'��3�ٍy�XEbi��G$<��;�?0�Ȇ��T�f�-b�8 ��!����@kL��d��
�&��+��� �͛�l:�u�C_�lծ[@���,�B���E]��&Б>dS��ayTK��#0e2�L�!��U���3�6p�� ��밲��6�Z�@4����E�B���5r�,ls��P�\��|$��1b4�����é'�����YU��茨�jZ��#��!������?i����I/��
�I�E ��8�I&K�朞�s�^A���Ĵ#01A�Z39@�}3���v�vVlB?1��.�\c��[�q�oӤ5�Ͷו���L�
p��j��������m����3+e* +Ny;5��)پf���rˢ�tsIh�����`����}f7����
�qo�=v���s9? ����C��X�֗�:G�*r�
�5�؃~<�Nȑ��J�򶾹�z��j�$�I� c<�_��R4�Q��g\�%�G C�L�H��}P��6�L�0
({Q�4G>ol�{�<��&�*㘞P��-yA������qr��i\'���Ж^%XW��F��� �l�Z�!��*���d'mE�w?WH2�����4P�_&Z4�3���@E��&1��� �b�Rה��̾������f\�i�k)�:��LUW{��ɻx�;m�.���u�R����e<U�ھgȒ:�+}��t����Ӷ� ���\K��N�a��-̍��MAgЎ�Gj��껗qߑo��B{�]l��sh�f�w]I�����FMPM��q�����an�B
�����X���;��������P���U��n�ERmw^зG��\��0�p��l�R�<��9���p�� 7wU`���������ȣ"���7�c������ZxvY����俰7�R�^$[���$�ԇ��t�{���g[6�O�<*ZKw�~���>���"A`b��)²4	e��s���@n���>�O�濾
|Mx
g�e�ߌ��d�"S������]h���U$�%8g�W�m��ޗF�b��p�bU�Gnr�IӴ����ƙ�ةt�zR#�]���x�:�Qnv$��9��-ȗZ|6v��:�U+VBZ4�O��5����'�>H��f6⫛��<:B��Ȯ�8*���ل��/A�&9��
B�b����&R$��c-���W���y@�]@�����sXT����|`~�t:|8>�<'�Vg���sT�Ѭ���P��S5
�������۹�L=u�3='��+�Xo�z�y����)R<�~��Gz���Ȝ]Y,�,B��^�QԚ �"����N�H^�(´��]ʛbp`�� e���e]�//�"WN���xʏ�K&�su���Ű�R-A�d�-[��-���e�U� H%a {�<���
�#�_�X�"TM����:�\@W^3E��B�w�Y�=驁�9AOWÉ�%�݃U��L���S\�<���G�`��Qs�.��������=�Wy��H{!�/Z�F;�_�Z���b��)|#�s�ȥ��s(,�x����w�~�������]1f�K�%����~3��4 �s�4>&z6l�?�>?�_�4��if��	��m��� �9:GBl�ikJ-f#!��`�gMlµ�V�b�-p��X33�>������:��h;�����`�N��Y��L��R��1:2>����r7$=��[�&p�+��vxQ��/�=Q����
�@�:�k(�D���A
�R�6�.zB;meӐ���(�
��14,-����g�ڂ(=�Un�ߤ�l�V�w��R���V��'N�� �B�A�H�-�� �<�8�|4�4!��e?�3~xDn�W�#3g�w{~��q�E���H�#X��L�#�}QRu�KBdl��ߏZ9��#ׯ�.����N	�ε�4����T��n���Y$XVsy���qPt|���B:MB�{�c ��B,�<�0f-`�Z�[SٱMO�l�Qƭ�_f�LF�n����8
rM:�l�J
�q֯ @̮���	��˳��0`aͤ�Xamt>���xp4�a3���V�v}_��w ������ꨫv�7�k���`dFF4�XlxVHYEB    f314    1b50�'��Y;�p��2b�\�OZ��0�`�b�6�u�b덬�rs�K�&��iVޝZ-�#i/ZC�j�v�r�T� ������Ǐ�7�IP*�6�e2���x#��aaq½W��3�%��g��M�]��$��N���{ ����	�N�d��6�bSSPO�*e�ZP��F��K�jG����� �'�/K��/$'��Ǯ�H���?�	�5�yoF%�|���5^$/N4��O�Ъ}�c�W����K'���I�n�Uw����p��Xd�W�aC��&vJ ��1�� �2_�B�(D��phӌv���]`;OV�
t� ϭ �k����J���
Ah'M��,�rx�N9�}͆.�7�b�����^����l[�*��[�G��~�6�f�|��I�9��n�~�����(�7�^v'�M^ߚ�0�����?�3 ��G�_n���&�S�o�W`���|Z9/��Jg�(ٳ�^B`���j�0��mނ� �+�����3�]:V}����ft����(���]Y�/�	XI�6�h�҉[��\[�^�4��{NR��?x6�g��(rv�sԽH�辚w�&�h]V�&`�Y�<������N�f��:�x�Ȓ�j>Q�oNZ9���*��:3C�@��a��0�ϕ!�J߀���ݬ�������+( H'��~�EΙ+�ddY�0U䃾�ќr�n��&X�Sh�/�y�-�@��V�x��a
�AkZ�j�	��.*dP�Q�t��|�[�D�'C�4Xy[��T���f!K">��|E}6�izfմ �� �Db�)�����W+5��8��>�[絏XNI�1͠�d��>]Ѥ�̝V4�=����$���J0���:!��җ}��n"��� �@
�v�GUH�精ow�7�}������ݥ��J�c�7�W?�?9���1q4)�z�6Ɂ;ƩBQ�Pٟ�장�p4F]ǐ�#+����G����,e�K���t݃���X̑Gʾ>��o�c�j��(9�!���)Ώ9ɦ�����;i��g����E����=��j@0���yf�Q���L��2��5*��������
^O�<��~�e�!	BW�0��<�{}l�1�kU���7�*_
�tM_TQ�ki�	S3aj����}�̠��*6��\�[3��)�d��_� ��FM����q6�7��L���Kkf�4#���p��}{��D҈?9���O�k6d���o�pƕT� `p��[�{q2�NP<�	��ntA��ot�Z�j��ޣys�R���ˇA��$D�a�F@M�Y�3?^�"l��ꍋ���)�:~<Q����s�˻t����$4C[��e�;ΒH�_\�G��;�T����X�l6���S�=�=��$����k?]BSc�OB�+M�8	M�y��Y�Ǣ7/��Y��\�`N��$���v�"�0AMfVG*�8���Z*[���	k�2��L2�i_��WI�z�U��
K��L�ܻ�L��0g��~��WO��oQ�������}�`�U;���h�L�����t��uL ��0=�7�#�1����^<�``NIRgʛF���mfC~c��L3��fRpp4Vy̱ w�>Qz�li�VF��Ȇ ��p^��V6��\U�g(��.%z�����6L`z>;EI|K���?U�5��#-�'*��7�.b��xn�,>�t1&&���;�%6��5�-J4���.�
ⰵ@��Z����՜�|���?�x~'�%���K�ſ�pi��2��`$7��Կ��֚�$X)��Wc
؃���
Y�p��z�����ƽ�{#�Z�����ߢ��0?��8�����o���Xg?��V:����E�*>�]7)J����,�U�6/p��>��"E{ƥ��tĆ�U��e�K��q_�]�I���;.�V�8��tP	��:�z�{�8�){3Xc3$�-����K���L@Ij`'��j����~�F�QT�]ُ��B����Z܂_�TN�-��|f/���˘��y�,?3����/�̳�f��-E����ǁ(���[2��&wZ���~p�Y�!��}v�zw�2��|i�5�wvt[<�Zc�`T�Qs!�)�����"g�h�AB�/;����,���t�6���A�]��w��%�<)�D�9�<��������Q�Jrߕ�T�@�)�7 ��n�J�s���$�M��e�nǘf+>��)�~���az������Oѻ��@?���1�a<ԄY	��b�)D�v�M�͂����W^��0m-q�˿��_n���{<]��R����2y!�sGQ���wFrq�Z������37����j9{=_6��,�^Y+�^����k�,|���@���:_�K�j-ԕ�<;�H�!�a���\jTqg�����{&S�����"iEZ;`yx�|s�,���
z���3`���[��Ac!Cu;��_���U����A�y�Qt�s��2��u,��V4���|Յ���]]~���@&.����
��3�ȑ�x����f�h{��[��k��mV��d6�>!��ɀ�܍M`�ּ���f��&h7~��q��&��児lݚv�-Bغ�ǆ��4�z�`���;\�����0Y��T���7�J{bj��ßF��<f-��S�"�� ��W��[x����������̇� %Kħ��������Ͽ۱�$�pU�N&�Q�}ޫ4ł��p(�,SI6��4iF��z�Q�A�o�,�#}I�3}Ne<�}�B2����bo��9�[�L��*{�r��� �٦O/������G
҆�R",�Jb����G"�8��"�3�O�Y��+�%�����}�E����0�}h$ ���!�wn2/`� �ޜ��j�o`I���(=��K��-�>�:��+UE���;iO���$��@��GRgݛgte����1�،l��waO���OC��������@;*#�"T��� �XaQ��ݷ�`||��<Xad'�"�J��׻�˸39�]K�:|��˵^�h~�r��0���G�,O�Y2�]7��rqT�m�B̨*��KwV��
������A�i�0׉��I�%�Ú<��V�u6\��v���}-��y��D<{e�tD�'/��i!%�1�1!��O`��f�$��H��sVWj>.ū�fE��;EP2z[L��H~�,ƛ�7Լ����[��r�A���owq�/��	�����^�9��������P�<EhQ;n��H&�e�/��Ih�o�j�6N��>���� �5����?1��V�H���!�k12+[����A�� �k����п�.>l�$J��Z����W����QW�E�{`��A� ��TAN�Ƈ<Z���[ލ�A���Խ�ǉ���4��wL=z��t�j#��wt_&����2ȷ8�h�QG|�[$�.�sسE}�*�w��ӥF�?3�}�d��������D�7%|!�.�"E���m�e��|$�	}j���Y��ɴ^�
�ٴ$�%뱝{�OF��7��uc(���:���"���VL�<��Ĉ"�X���n��#I��A������ �#�Q^�۸)�1��"0���\��� ;z��Z/�XA)	m���s�@FY ������ �\�Պ`}���bMz�1�/ �w��l%d�B�\h�)˪�r;���!�`]l�,����M,U�z�|���ڟS~�l���т\y|�y��V�w��-�[u���38�&VyW�?�w�L称eq���Z&f;�&ųPJ�-�\��JMel0Gձ�$����:8�IL-!���v�+��J��9ט��0Ιg
��=Q�!7�L��y�\]-%���}��PG��4�	^�©Q	B��PH��̪���餢ډ���h�A����edR���xI�i�F;ީNr+�y5���S:bn���pz���-=��}�uu����T��O�D�`�q��KnZ���^�0v�����Refb>�ұ��>����GҞ,y�O_�oS-΢�x?� ���Cx����nϋ5���ݽq�έN�����%�i+�|R�*^�p��Y�����0'�c|���h��4�ɶ�4A)E���������D&������R=���|v.��������ʖI��0X�zj�#4=,�F Â��m�$�;�NJf�}�B<aDG�m���%��#y�:��Lgv"3=R�Pw���=�����������6�TQ��z��65~�Y��h��QjK(�/f�	�qP�����<����4=�ݚ��o�;w���8Ÿ��]}@��0�/-bvp!��2�شæsߣ��
ٔu"�0v�0�$��vd,jn\��#�6�� ����8C�ҋ�3�s�����m�,d|S�B�=)�w=�I�Vx��ͻ�%(J�O�Jz�&�s�4|��B1� ̥��8��k��т��4��{����J����#�ޙ��m���my���'�
��A�<g��uNA�e}_Αd�Ӿ�z?L@q1�[]���r�Y�	��O���^/��sx*�T��K%I��DM !�pg����Q�n����7��O�5;�d���h�*q5�Мw"�I{!�L0�R�*�Y��;���}�̻��F��V����'(*6UB �~�����жe��Ǟ �F{� ��x�a��A�ԝ2��9�/uQ	*k/�|�8���� 8D���Z��,$uW������`�FP��n
�Td���
�ob�)�M�n������S��=�	�R���:��%`\6��ě���\ht_Jo�Y�%����,ki"���C5W�p�7/��W'Ί��x9�PUp�P��mԬ� �tt<��J=JO�ݪ=q�8E,8	����;x 9|�%)�C�0�[�q�ʭl���� �IT?��0�@*�����C�09M�
�bGD眩��;��a_������*G�Oo�=������W6��`�a1 R��HѠ��x];M��v����\$���aDK��B��<��X���8��q��Q�y7��ίr=,햨�(��z��CA��M�X[#�<�����騄l&��*��\Q|��� �}�	>�{��L���)�A�d k���T��g�m��Gذj�z�3��VK�'�0���wM'b��ݱPޝIx�T��gD��:2U'���˛L�#�]՞T��Nz�<E9y%�Y/"f�yβ�+>D��s����	��M����c4��F��qJ\�7.�����aK��BL-:����ǐo�Ѫ{R%��X,�]l߹����S~��׌m�� 0�j�8}KQO~ut��ݺ���U�RZ6�j�=� �3����x��SүTH8��"�VSs�+���&��1��2m��~&&�7�1�f~��W�\�� x�?�v5kQ[�m�7�̓����	��6�"��{��J˝��.��kc���u�@<����]�����m���:)���5O�d������x_7WG U��m��@
�l���͞��<2@�����4  <L�c
�_E���*0J���=X��K��}�<}[�fx�0��2[��C��G��&��}#K��N��5nԗ%>S�)&��0�?��Vf�;G�����҆�EB�^�f��6��fx�g�B̛�e?�yv���?k�r��&"����rE+s�Yr[F�jrF�jwL?rv.uE�kBW��5���ϣ��!�X����E�V���E.zHr�nh����:!�n��	,�Xtv��p��y2keX/0N�G0xZC�=i��o1H[XeX�x�2[�yϭ�w���m��Z�l�/�SK�_t3�6���s&3��&Y%j,���-Wv�R.�9D�O<$鮈LהF�#�gn.d�]�mξ����a�ĭ�o��|�|"il8( ��;�C�է!��ߧg+�:s�h6�-EN:׶li��S;N�Z>��U��;����U}m�=���D���Bj;�D@���We!����v��,=
3݆3aȰ]*0!�)�l_&�V%��hc�� ka Q�a�u�a�(C�p�>���ȓ����u,�>����˄�����R����f�x�~&�h�)�}���q�g^9B#pߎiF��g�:Ԕn2��=Ə*<�B�'Ig;r��oR�኱Hl�f,Q��<���7X���\������<&/�_��Iq�6���J7D �d�ݜPY����w�J0��Qej���ݱS�B��4���g�b���e����:�f�3��!�c~��"�43�3��1���b�����Z3�@ �.�����Y���Y����G����w�.�ȝq&	�R����_Go��fK�n�f[��eѷÕHk��"�2�P�@����p�B��1*?Z�Ҋ���px،/��_̩7�܆���=Wm�F�2���ע%�ot�n|�D��. ���E�>�MYr��j}[����
j#�5�M*����F:5�	��}}�w�w�ф	�,A���R�)m���������*Tk0b��l?�)B%Re�N݆��d�U՘��W���>θ�F4���|���d���ﾠ�S�ZZZ���bAys9��R�������������+_����C|3,�[�_/���߲���f��LS��'�[^�?4�RX�ɓ�F��	�Ķ!��v�X�v"^�Z��*`�9/J�QJ
vhm���	M�\|FK8;r�j!�%8�a�]��.j�0{j�h	�c��ƌvX"�M��Yf��K�"�6�)�N�����م�z&û���Bg����vCx�'$V?�φ�F�{^�T9�\�����5������x�Ѵ@,��"�5�-kΣTWz\'e�6b)�� ��]