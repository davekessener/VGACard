XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Hm�D�	l�AU�Gz|��ڀ9CAj[�q�O>����Zϐ:B멩�zL|���獉����߄Z�����p��Z[F,�N����o�dr�{��9�66 &/��3��nЌ�L.��f� �Y,�1	9T}J_��������g/23���D��0z���%F����`�Z��ۗ@r���w���x|]	g���)W!�	��@<��	d矬@g=��!yش�1���
t�g'|�X'� ;{����#���'^]X??{
 C=���)��X�����/��X�.Zy�5�"C����jW���!���gHEМ�P�*�$ٰ$�Fob x�p�Vk�mϊas�U-�T@�9tCa���Q��u�fg�b���l%1n����e	"`^��8\2X�N��������ߝt2����A��|<�VGGQ�Qpo��l�T��v����x7`<�zd�Y��s7\�����ؘ�s[@�b����Wռ��.���8���.��_�vi~�,�'@�5�9�t�$����[lrOT��Z��>�(��[���x�lLʳbad	�VM��j[�����R8���gd�c���a'���w?|�p7�8�͵^�Ul�͖ԥ�X<�衩�,,�I\�'�ѭ�)3[�A�U���6���!�'�(���a�1���C�B�z��
��T퉄�_o("�"��)�Q����ڜԢFr|>1X�>���N^!w�JW �(�ċy��<[V�e�n�� �2f��#�ƻ�o�C��XlxVHYEB    4089     e40=�!�ӕ��@����9�x���\�*�� P��/k����{���vb�qĆ� �:�W ���$;W�����i���)2U	U�"y�@���٠!���a3��!�ƒ^ҋ���?F.PZ����OD��d���UT6���d���t7�X��8Q�a����	f���+�_R��e�^���(:R[
�ZQ9�Јh��Kj�f"�䗿�]��P	.��	v�7�L�.H��|ʷܱ��C�MNS��0 ױ��u� 8�S�m��T�K�L��&}d^XS��!��V���1�m<W�'���5�m����W8��D��<��A�N�"�u�쮹#f��G�3h��n�����En ��)�_��9�
�3%ʩPf�"�u���a��J�ۚ��]����V��a31w���[':�K�^;]}6���3��KN�/��]_O���IY������hs/N:W/�#��Ù�����~�Ю8��>;�w!G�k�������:�<�!
��.�tp����B�*��+A��򱐬h2�����&.��6�\(s�u�!=ƶ�������(�X��F�� Y^yϽ	�e��z��J����u7�Y����ӓ����P��A{�;��B��je��1USB��5q��kK�,�x�g��̱�Ke��[$��We������yN�m2')Φ���N�C?�i�Lg��>8���v��yP�!Bk�%�b�PÄpV��Bn�w�����c1:�J:|��@b4�s;��E٭?���9��:��a���Z��i`�]����6�C�j��M#�AX�H �rZ�s"�kUӱb'~��Vs�e��Z�86��W�f r���M��}fb���Ӭ��QZ�!&�B#�vOz����3t��n��~\ D�f��e��@�l����Y#�Q���.�	�z�>L�?�4ڽ�!�X��~	�S��K���Luk#�k�.p}������qt�Sξ��c$8:��q�kkzXy3HE�L�:�,*{{HAi))`J���/&5	�`��z-�rn��т���߂<z�ݻ���6�71L�b+b��݁��?��M���P�o�sY<�@h�� �d)s@S���_�*�zR���qG�E�䨀��U�1����Y%_`m�����!��'��"����è�p�d���\e���K��!f����f�'i�G�2b6�Ï�\�\���s�����Y�TI�S�d��6?Y�|Ǜ���ձu�� [��y�����~����Y:��uL�m��e����R������E�H�%д�O��&�[�=�����P����+��	�:�^�����H<�D�A�F.�ܫ/K�GvVq���+7�%E�������Y%Ww�������iv�S��&<����8}ST|��9���á�^�<mk9�bq�;1hsQ�m��j�8���TO@w�p^�47�g�̢����e}��<�6���@�,"�&��w��������˫m�k�LV ��0�]d��KܹG��&}=���G	�v=���3��O�/�(������)�3����4W[�%�`��V��~�!Ĺ����f�ހ��-#�}�2 U��C���5H�����d�6��{�N�.��,�
g�f�B.���p�+��� �X�J>)u|��Kus�*i�.���CU��h��	d���%VZ�5����P+�K�#�4A��?��^]�3����m��&',n4�����>�9�������5˖�TPȼ��w�����Ȕ�b\��]�LR�o�_��֘�8�}$�� m�r��O|�C�P¬Ƹ�*��6�% \��j�۬*���-��&9�䣱m��������q�J�.>�<&*���8s*��LP����&���T�S����ǽ�����L��}��c;� 8�"�*SM'>#=����/�#=��>ǋ_�cgnwB;�~f�m��5S����{G�U����\5��4v�I��⦇~vL�uy#���A��~����m!Y�G(" ���yy2F�%J���# wO�ԑi��)�`ʫ��RT֭-����f��0�5_F��\���}3��j��6f�}�YXշ��azխfnh^z1z�lw�8ʪ(��Z�4��m-�6�e�'!�y�5��w-�&	�e�280M�[_~kq��2���9�;�,���[Rw5�|�K%`1�Z��95?Q�.[ӯ*|�Y0[�wcO�@�K�𚰣+hm��A2�}������䚃q�7���J�FO�	�6(41y�V�Ӣ�h�,j�SM��,���(0�W����x�+�Ă�]���){�w[��*�c!��aO#��C��*/�a=�-�G��Z��4�:�-�B���V��/����,2Or�a���/&�eB�<�4$p+��#b��̳+;瞴���c{�&�gw�B��H��u�V�r�`v��1�Q���Su�L+��l�+.���ct�0�G��������я���che|k���䷓��H&}���gMP�)l�l����/~�^)�7��Y�xR���7��l+�)�`�$��j����Z�y�~y-�74�ض��5rʩ 14q�J�L}��eQڢ62�Xn4�6�� {Xm��
�{BD�ڹ���и�
����F����6�0�O%	��`��v1��rD���A
ִqߏ��5�8��b������kK��#�H!�O��ֱI�9$6;��!%/����3�}���$�v����m�E*#e;��T{���p�S4?��7��v���)4w��u�	=B�H��O��C�8�^1U������Q���G���f��Cq��|��w�!��}MU�C�ƀ��1\	!��<]��M��Cm���霮΅���2vGة��rl��-����h#g�GZS47+�
��_�R���=x��^��A�i����r��]iM/S�l��o=�o��{�����a��lL��c%�*C�����|i��i��	�w����Z�]��
j:cpB�6���A�yg�m�I�u'��Y-5�I%?8���:�ic�Ϳ�ٍ�1�cB5��1l͖�zDpN#K� ��x�!b�W
kG'���n����
BD?J ���q��g��7g��N<Q����S���]���ԶϜ�i���;��O���qH�L7&�o㷫&)�2�w�C=ՁPX���(�U�W��+�����8���ۃ{�Pu�x�񾙷��iGvp/���CTxs�#B���~�����Yc�p�$'_Z|0���a�O�+��?dR�v�a��Q^����9m�9�y��,ÎW�Y؎H�A�꽂D��! ��Z��Lv�+����Z�}����g�Iu��� ;4 �x ��Z$+���-�Ki��.yۉ;B^����J�#���R24=U�J�Vi's舷0j�w�fzTY�G�n�N�i7���_����@`�C������BvR4IS_>áM[�i"��� B��"�@Ĵ�H��O	�<_仫��F�-�<
�����4�/��\�|��KQ�I��r��Vj&,U坅���uG&s��E3稥 '{�^2�~�3�r@�1Х|F��s��?�S�H.O���S91��˴Z���G