XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}�m1�?��(U�,����u���@�IhW�[��d�qΉ�$�(�J	R�3�Ƽ���,َ|�U^E��\K�j�[6�n�ob�JEd�Q��p?��y�k7�;�ƨ�+��j|����M��ʎ�|,X"9<tb�����q̒wXg�@ ��� ٷT���=���e!ҕ�W�2������s!�,)��%ζ�m�h%��=� l��[���D9N�%|k(���+/hS6�V||Z���HX[$0/-��h�������@y�D 2���I�6���&�1��[a5�/��y��\���[��k����5��צ���x˥Ћ�N�Q� ?�'؃p����6��9�}�P݉��n����j��Ǡ�L0ny�y]��-{oպ�	���P����W$����gM�G,s�eoeߛ�.������vs��;up��b�(X�"�+�7��An�/ؼ:"Y�����B�M/�m&(���p� /&�-HA�}3�ά�٭�dڲ�q��h��bP5C^X�l�yf-��Te�%��<;��)���|n�z�����l)u��'�:8E�l�<�����eۛ{�^)�H��NKC?�i��p+���&���u\g�D�@"
ٞ)3����(5ر�~��^�-���yok2�X�&V�9�e}Vn$�N+����s�O�a��{�ǚ����]�u��5rM�b�R�SB�]|D}�4T��f�Y~���h �v�'��]kW�Y�ȼ����]�"9)采)�vQY�9���ϠXlxVHYEB    fa00    28c0ؤl y��!����q(F� N�


����BCf.xC�Y�"Uʩf[�U`���zr���H��f|�U�ԶD M�?��-�]�l��c�ť����5�:��1u����n���O;�v �%��o:/��j��n�W�
k腁�M-�X"5��b��HC�`��g�/�[���笙k�'@���'�zhd��<���m���U��]U�����d�L`k� ���Ƨۜ��m�K$�D6}z)����i���[��t��.�;��jD��J�ɺ|�i�8
�ߏ��V�2���&��Mir��X�����5���úO?p^����!A�"�̩
ܒ�����̣|�LIӹ��
�53F{�ss͝�8����x����Y%���	Ĳw��:��7���9*�4�ʯ���iQ`q��'��9'��-�ͷ8�\:��E�e��j�/[3���I�%�ij�帋f���K^	zq%�qx��/��o܋ƳU�{�:߮ �V�x��Y�&�����O3���;Ylo��ۧ��(��ȳ�}=�I�.C@�x��t�m;��I�Y�*I|'�W���֓����Ϣ���9�d�g��!�����!���!~1��K,���S��7k<?��
[׷�k��X�3#moC)�c$e����~0���-���Pwe�N��K[-,���2��y��&��%F�ߨ�A�����>l�������wsݞ6��w�Z��q�D�-.�Oߔ����������ƺ�C��B�/)9��_���9ۨ��W"�%��ge�m�0G�Yi�ԥw`2�뜳nrnd'�2OC��-�V5!����)/v9���A���(B��$hoA�����nj( l[\�u{����L�y���#/����<��{��ftͻ��VgO�?���_pM�&��8��:ږ�?~\@�y�@2T�w,[6�j��y#MVW1fE�!$ �x��g8�C�)%˺qb>���ԅ���)��0�Y-l�@��'�\�5�
`K���\�P@�t ���ؑu�����{�;�Gt��[]na����OQN5�NL��W�%�K�k�`����&����K��R���~�ե�������_�Xҹ,�1!�z�x����5��f��8!߲��̇�xu�|1F~��+}%��TN��8Tro+��)JN�ldn(�N0.��o���\�g.�L���wD[�ӂ^���_�ۥNC��g* �C�P�f�n����X1�1H�2�B��4�1�<�1^.�B��#v�dHP'!k6kh�m6Ы�]~7��ħ�/��倂NH4ŽN�Kt��lTVpΥ����A3QWG\��l�f�i'�˿k�U��b� ��4��H� �!���ǣ�(-0�U�]/��dA��l�2۴���p��i!:k۸�Eh�#����_��	��h����w�!��2�p��iN��R�4#N7&���n[.@�Rە/�:�7�)�ϕ���6 k�#�j}�����t1 7���c�����ڹU�Y٩ R����d���r-�ܱy�o"BZ.0 �V�Z�kZS���W�Z��l��/1�����#�֩�t1�R݅s���_hJ襾�Hz�� 8`c_&��Uu�j�	'�� ��7��X#�e+Aq�����P��3�(������`��3�r�*߻O��?��M�W��׌���|S����:��$Ð'Ƚ��J��F�Ehe,eE"!�U�Hk��F���ӞU~�_<�e�u���Gu�.�����s�@����~�x\�A��q�J�x%o����Y��w��ݘ@�IO�Ƙ�`���A�xa�O�C�r�h��Ҝ�n��Z���G�қ�pv�9с����$(��*����MC8NY;.�r�[m�	�2]'�	KG�)�XP���0Y(^� �z�z�;Y*�����Ѳ%�
������&�¬H���/�7k����~0i T�2
���1�^ҹ�gg^�a.����ۭD����whj�:�ء�_���Y�/7�B_Ǽ݄J� `���gs(�J�o,�XY=!oe�{�meK0��:�B��Q��k*X�Y���� �*�r��H�
��[4�1�����ܾ�h��O]x�9����A����-���w�7����Cqծ���JA��[%_�j��
��֧?5�\k߰���h](B8�J�^ǐ��U��k��/����nrvYr�_:e��]����G ���7ٿP��
�^���dG\lE�!���̔j�5��E��X��M��P���be�W�iĄ}��%��1�����e��P�*r��q�)nrW
8G�m��է���o|���X�q�A��������Gz8�� Y~J=T�zVp�G���I�(|S��нdY�I6��Z����~�8�za+�36��]nE���쏵{o�������V�T����)��bS�˺̕���3!,���]ud�0%��N��Q�d�/I�m�p�i��gX���k8*}�������*��Ԫ�4eG~�~�M��M��Y>��wtxȗ���M:�N��}��+�B��4E�wp*���9�%4:���)��h���HJm:5Ae�9�@"���\�s�;�$��;٣��
�'R�vp�
^��{d5�����d���W��RWfȞe5͋%K!�D����^%L�������qm�YO�b	S��=�@n*{�!�/�ef�!��nwr���.@�(�3/"�J��la�Y�#��å��v�Ծ�}��IH1�)G!�m�ǽ72]:N���̅&iC5"3ډ�>�;Qx�ӯz���eE\2�B�����͸G� v��H�=�N�I�_CѬ6��%����<=/� �8�V(*2�'O��5�L�!φ?���Ʃ�𭀠S�&����/��-�b�
ysy���Z@�f�O�}��,��D�r,E�%�2��HI� .���řU����s-㏆U��A9t�Q�
��K�1���`6�T1���KZ@�R\�;�[H#�]��P<a��Φҿ��y���[����-��]Y��bT�$��'m*�˙�Y	x������<$��̗R\N W��0F���{(��<�g~?�i�ʵ�y�^?�
����!]��U����W��(JE&��	i�֪��X����ln_S�b	�$��G'Q:ԁ���0r�[[B���*� R��1Ä�If�vv9�Z�����-�
�`�ߦ0#�,s�Bw�НMZ�O<[�`�;~�j>�ۡ���+р�I�d`}�m��W�Xt�~0�X#0Ԍ��ȼ�g/3�GĔ7�h��	=!��og����L��wi^zY;�w0"tٲ��D^��iN�p)<o�d�B��0�}��(R\5���hX�ꊧ�d��/�^��=U-\�;��U�4��a��jHO$�e�m�1@���G�����둪;��#�錫+�������3��n%����L!םo�Qzؕ1N��
N��s(�긌^1F¼���.��^��yƽe�<Wj��i$�ˈ�Q4��K �6F��ؑqw����%V����e��V�(����/%�v>�YKSЗ��#���SK`���Xr��j
�z>F!*h7~�R�HZ�A2�o1�'�n�aB*�ⱉj0@����"�������_K��ơ���D�"sٛ�PMQ��d{�H����Gl�m���Eq«���;��Do��n���x�U��fV�'m�%�</&δ�=�;é�����9�aJ�Br(��4%i������I��u�C絩�:�^��y.pO%�wt%5�3�J�T������󄕊I�E����_,��V�v��	c��0�����%r~5jcR2�y&����7�e����~Άrɷ�r�G�-��$�+��Q8E�����Y�KzL}��w⢺��Z��x����箥?a~g��}�!iP6 ��p�nd��)�+��&�j�Dz��#o��O	�����gު�Y�:��Sgx�#���� ����"Ր�j,��nd�hN���v5¬&�x�΢����������D�"��&[�iCJu� w|_\����_4��P�`t��]��RTe��hPx���?P�>�M�B�g�.U��#�C�0�l�N|jX�VU
�Jw��v;a_#���Ka���Z��S������쩽hr�2'�kW����ie������i˟�u��;��������/Ϝ]q9����>4�Qy���a��Ve,l>W���J��m$�êt�Dg�W�b��.�YW�ܛ�z�e�)E��F�e��ߝpZ��/
-;�Җ��^O��� o9�?��FR~O(g�"�v�6�߁K$.����Ȫ�����>h�"�?�n�&�ύ��g'���<�C"�߾Z��R�����e��7��U�����S 7#e����.�t��B�� cך�cdN��o	}⻷㶓�8�gj�̯А-�i����;G�a1�6T�{�`v,zi�{kM�m,@��v܂ۨ!A���r8�^1
	d������@�ϥ��/��k�Pggڸ6G�Ӫ"�D;=�nL��>"�ތEռ�y���������A�{5�y�����y�	y39_�/���/u�.@H>Ӈ8��v���JR6�3�2.�x���ɟ(��D����_�T�tL�"�8��h��/$4m��6����w֮�+�3ir�}O��#�]On���D����Wq���K�t`� u3�M�'{��\,}(b�[���#�����4���i5��@z	�����I���$~kߥS��kw�n�a��.�FC�����]C�D˕D������G�.e���jN��S!|�����!��p���<bg,&a1p2<@6�C�.H6NF�TO��w���P˴���*e�x!#�'XM��P�!��
�ݪ�{���.I�5_�0O�����5ݪv�P�G���]+�r����z.9&Ŏ� ׊�Q������/�ʦސ�uWB�^��r�ibkg#T B��RڧPВ�B'5�_1g���)����>H����^�9�<����e�2���#hE�sM֖�+D�*6�86��U�q�U��f�'F���|�$��w5��:���@P.�ޒ�*i���;<�����3��hˏ9b��R���f�ADE��`�pe�F��	�n��%,�����t��R�԰(��Nas��0��c��"p7ElN�Z�&��N���N}�8I�_����>�Y 7��-��{К�EDOk9�F�P �}8Vp_FRu=ge�	4'j���ˉ*��9�OBc�ؖO�/�h�_Ƹ���HE��q����$��9��r!$�Bxc�*� 0��G�vEOrs���Z���b採�!����ޅ{�2�Na�<۬@��;ԓp�w�����򔍁�]'c��۰q�F�~,��q��^��i��J�FY�(�b��Μi�<��`���-�GK4�y݁�W���ꑀ��|�s��w࣎�}�jL�6�?��'���<;e���?2)$�v��aCQ��)<�
��;�4�C*4��� ������"�M���Kdy>Gh�JjA�'�w���YGN�=7�}���k`XKP��ऒS���|	!k�3�]:@�5>rwi��@Cn�A8�W��c&�ČC�%Q�R�z*Ҏ����H5��m�i�kp���Ά\��Nɖ�$o�{�k��Ge��A��QgEl�T,= ��5O���6.��&�����Y/�OR�u��ȇ����k�`�SEnw'$��r$0�N��e�:Gk��iU�Uo|�vw{a�������i�1����Ô�&ka*LE��,��f-3���Y�� ��y0��b�y���zH�����5R/�s�Y7��i���7�;s�5����̀<���F��6'�#��X�+�������3@y�V�0� �%1 ^�Lb|d��p�|�t�aEc$���s���[�5�v�m�fLj�w��|�=J*)]��,R��O���t�W�g��|;����5�\ĊJ�~~�@(H��l!��>5�ڂ�`�Fe'�ȌJ��s�pD3�1a%FqP��u�e:Q���D9e`	�5Hj��&̞g�;-H�9��W��q�eO>#�1���X���������p�>�\� ��a|:�Fe���}�ߥZ��D6Dt ����}�o�Ё?�6�K������!���8"����$o�K[�R�Sf��M�h��u��7�:\码&	��i�_fβA���_�Q����:��Ef��)�`�ƕ�����dϋǤ��%�Ʌ��ɻ)'�(sԍ�0���j�7�(�I�Cs�g��������ڻxZ��[,4v%����:���z��x�"�
�����������>ׯ'�N��TU��� <��7��$;Ǿo�VK��Gc���5����SۀB���k�,{o	`��OŢ��T���F��¶m���jO �p<��W������$�
��, �Y���s��D������gn�/���U����F��`�W'����i�F��Wz�[7ȝu��g>���?��KDz~�GB���Y�Ю9�����Q�Zr��7�:�^�����W!�L��]:j��M�)�3l��G�\A\��ot�,�47��8��!j�\3���u�$}^Pi7`�<P�u�u��:kã���w;J��b�j�q{���<;$֜%����3 ���z�Aҕ� q о���)��a�5�P��q��9L�%�mDOK`
���0�}���ϒ�#��^/$19ø�����:����q=MF4�9C���&I�F��FN\6�G��iD��T���6x	!m(�O������%����ܖf�&J͵cȸ�ffl�f������r��V�_�dY�֢h�����F���B6��q�i��e]<~+5첓��0��!����=Q���0�P�t���r�O(�M���e������� K$�=�TĎ�"��/��)�G�&����z-�����"�+s� :��:�5��ߜ���|>�L��(7��� Vn*X�'E�ڥ.p��tA*�\���kD��S&\-�*����e���x�Y9y������ӉR�߫M�����_�bf�UFXΧ����o��T��᜛���^�zAʅT�J�r
��Z�_A)䆛-_�xj��,��Õս�-�7F'��]�g����ὔ�g~��i��=Gʉ��.���*��K��]��Y�,���	�]zD����Nb���8nI�)�����`�%a�D��8(�@.n��7
og�	IF�a^���K+�/�BA�b�ROD��6::m��5Fl������%�)�W�fVS�^�����L���iZy���0�P�R\��a��YEI@�ޔ� ڞήw7x�,.���*��A�)�5�9Pi���"Z�����Z6<VϿ:6���CX�#^"! G�r���k�&q��B�V��?���ϴ��)�x��?a$�:)J�~�]����v(��M}A����D�TR�c��c�Wc��1���43�171��<�~27��o�k/}�+�քJ��)�/����i��Q7�CY�H��9n��#�(L�Z[8޳/O�acw��Ug&�Z���")!�/Y�ߙ���ńݣ��G�"պuv��t��E����6���/�9^�'��v��(���f��O)��Z?�]Ox�r��\�%�ίm�V��C��p|��ם��OP��+��U6�[uꤿpX��4��V�IhńE8]�i��'n.�FY�{
����dF���I�;Ϯ�0�$F�6.�p�%�aL��;���䍳�A��nC��U�����雏iiĆ���=�"�ͼ�8#����,�����h8M<G�#0����I\���t���XӴ��r��ko�6]&+6~�p���3��7Ys&̡N�b����<��->!�njK�G~�J�:�G=hy��Ci����Yϧ%*�[o'�Ժ����)�9�F�S���H
Jl��������evmU���,#)^���y�n@ѾJ��Z�eD��#�p(�/��(����B�(�]Rߡ7�[sF:,h�>��|�:ϩXu>�꺙�<�	�����Ȼ�yF�/9kX��z���k����#a^��\�L)�[��x�G�jf��?/�ar?������!f�̏�֝�n��͙���Ҝ�����@����:�b�V�tpXcr���E�� Vt9IA���@8 l���9)'�S,����
\��\���~�XR�����C8��x�6"[��|�r�0�P�iحG�Υ[,?��g?#�,���:�C���
�T�
T-�7R�d����y;'��NӋnm���ՑGJ�д��� P|��+㜍��w�F���H�K���>����~��ʜ~DW/��x1���c��s��a�đ�3Rl��v߸�K8��vDQ�V��JI���Gm�%|�6�U������ �}�1}�v�c&B�vC�����i$G��١��wp5?�8�Z�ѱ��G��� �I��y�K �7����D İ�;�P%�A��z}��v� !��=/LRz�F���Q����\�2�|K�/�=���9t���?�Ջ���� c�(���r�ЈE�?�ˆh�u25�f[Ɵ��k~0�~�7k�Do��~B�[�*�
�Bܿu�d���ƛ Y���~�VJ��XJr*�]��/`юI%������d�9�=�A54R����/�A`��ޭ�W&�$�@��{ˈ��a)�k6�_+<��+s���|h���ず�3	���g��O�4�q�5�f?0����͔t)]�:$�ձ�l�x�,g�[G��g��S8r2때9���ڕqF�����1h�3�=w���T2&=�j��P2��$��e,B@�ۛ�� ���_�,$��!��z ���g��&X#ض�p�t��C]Z�So2'��h�@4���]B�e\{��E�q_�nW�����Vb��2\�+�����ؘ�������>�iB�4W� T�
k�KOЃ�)ȓ'%=]�j�E�9f���K�"�3A��Wڢ���0{���f��5�fL����KR{���^��zI�X��~�������9E=-R,��n�V�rW��W��GI���LoJl�u��,4j��❦";��T�g��F�Ar����]آb��""�_|������T4>z�֙�oy�� -�%��:Y�8Dݱ��2���g��O��]�N��-�f�Z����%7����5�u.N[^ ?�g�_;��-�����~1�	���D=�2���nS��H?���8�.�:�t�պ��!f
"�V>�2h `���g⣧�P��wl���'�K�����R�?�t�8��}��=ݓX]fF��=>��ؠ.�.%��!}���j��Cr6��v\?�ѩnX�� �Y�����C�?�x��}��oFOY�<��g����*<|�q��1��4B�!e]�7D����U߿����M�J��k~i�dךCc������*V�]��n�`wBJ�*ސ$j�
q�y݌�(��[j������Nj`0�\['��箶d�Z����ӆ�n~���$5�m@xU⚷�-�n]��?��=	vq��*d���"�����v>�T�<ۢ$JaTϋ�R�<��W9�^�YF�]"�3�a�:I��۪��E0�{	 �tqH|�K���Dҵ��7�`M1�A��B6�]�=���
s��#��tb�����ġׂLg�s���i<��B���a��A��p]�x�:��g����䗰H�vgx��B�tD�NL	C�*�� ��t}��1��=�̐IZ�N��W�v��!]t�ʡH*m�#0�;cu1�|�N{:�9K5�*�?yR�2"� �{��.WC@v�W}�Uჟ@*����-�yy/�~��`���P~�CV�4��i������ӕ3�/�s�i�cDp��-;5��B4X�iF����x2рYǾG����T����x� �`�9�[����xm[� ڭ�	:�^�~�`b����Ɋ\0���O/t��B�1��|��|>-OHY�~x�8����0d���l�\��w�F�/�
��Z3���P�5�H�N9�]���Q��d��/��
�΃�G�{�_G����ܭ
��6����{I�[X�;�̛�?�7�s�1	��f�C^kQ��y4��K�TUZ�V����D�ӌjib������1�Ö3\�K0lOg�ԝ;Vg@=O�J���2:TF��g�T��\�Z#��}�IɊ:w5��R'����6���w���FW��0�>XAIG��8~�G8XlxVHYEB     896     280�.up(QS��шe�ip�m�N�DEfH|-}6�.pMj�M2�!�7W}����)�}��56H�Q.+/�XI��f���QBv�]T�լPX^tC�V+��:�T����mD�Dz�Me�%H�g�+�B��:�ƗhY��f+�C(E��4�s|nF?���gV�٪��d ���rnN�}�?Ag�|�%�1pԆLS@�6��A*N�ܠ=;[vg���]"��o�37JA�yjp�M XW��.�S`~�S;+�K���-�-������y�[��� ,�xi ����2����?/���AZ�wZ��ީ{��#�/d�"Bw��;߉nt�Q^Ev)[�Ti�J�V�E^I,!���(5��wr�uW��P��	�����N1Q�1 ���ݵ2���M��GT�g�k�'����nk�_�\!��Q��F,2�C�~��:�{v�#�A"�����4-Z]O�����6�$����.w͜�J���޽������''�K{a��CS'�G���	�_�8 �#��r�F�Au����E	��^g9Qb�>r	f�mWJ(�s8��[	��'?A��xf7�.� NDH����J��#
�(���ն#�W��8E�r�6�z�K=0���\��b���Iiɿ